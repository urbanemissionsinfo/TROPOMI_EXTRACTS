netcdf S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919 {

// global attributes:
		:Conventions = "CF-1.7" ;
		:institution = "KNMI" ;
		:source = "Sentinel 5 precursor, TROPOMI, space-borne remote sensing, L2" ;
		:history = "2024-01-24 07:22:46 f_s5pops tropnll2dp /mnt/data1/storage_nrt/cache_nrt/WORKING-666967739/JobOrder.666966421.xml" ;
		:summary = "TROPOMI/S5P NO2 5-minute L2 Swath 5.5x3.5km" ;
		:tracking_id = "84bfaecb-7086-4b7e-9dbf-54daeec84ada" ;
		:id = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919" ;
		:time_reference = "2024-01-24T00:00:00Z" ;
		:time_reference_days_since_1950 = 27051 ;
		:time_reference_julian_day = 2460333.5 ;
		:time_reference_seconds_since_1970 = 1706054400LL ;
		:time_coverage_start = "2024-01-24T06:39:07Z" ;
		:time_coverage_end = "2024-01-24T06:44:18Z" ;
		:time_coverage_duration = "PT311.633S" ;
		:time_coverage_resolution = "PT0.840S" ;
		:orbit = 32544 ;
		:references = "https://sentinels.copernicus.eu/web/sentinel/technical-guides/sentinel-5p/products-algorithms; http://www.tropomi.eu/data-products/nitrogen-dioxide" ;
		:processor_version = "2.6.0" ;
		:keywords_vocabulary = "AGU index terms, http://publications.agu.org/author-resource-center/index-terms/" ;
		:keywords = "0345 Pollution, Urban and Regional; 0365 Troposphere, Composition and Chemistry; 0368 Troposphere, Constituent Transport and Chemistry; 3360 Remote Sensing; 3363 Stratospheric Dynamics" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast Metadata Conventions Standard Name Table (v29, 08 July 2015), http://cfconventions.org/standard-names.html" ;
		:naming_authority = "nl.knmi" ;
		:cdm_data_type = "Swath" ;
		:date_created = "2024-01-24T07:20:29Z" ;
		:creator_name = "The Sentinel 5 Precursor TROPOMI Level 2 products are developed with funding from the European Space Agency (ESA), the Netherlands Space Office (NSO), the Belgian Science Policy Office, the German Aerospace Center (DLR) and the Bayerisches Staatsministerium für Wirtschaft und Medien, Energie und Technologie (StMWi)." ;
		:creator_url = "https://sentinels.copernicus.eu/web/sentinel/missions/sentinel-5p" ;
		:creator_email = "EOSupport@Copernicus.esa.int" ;
		:project = "Sentinel 5 precursor/TROPOMI" ;
		:geospatial_lat_min = 32.02938f ;
		:geospatial_lat_max = 56.08662f ;
		:geospatial_lon_min = 71.52991f ;
		:geospatial_lon_max = 111.3999f ;
		:license = "No conditions apply" ;
		:platform = "S5P" ;
		:sensor = "TROPOMI" ;
		:spatial_resolution = "5.5x3.5 km2" ;
		:cpp_compiler_version = "g++ (GCC) 4.8.5 20150623 (Red Hat 4.8.5-44)" ;
		:cpp_compiler_flags = "-g -O2 -fPIC -std=c++11 -W -Wall -Wno-ignored-qualifiers -Wno-write-strings -Wno-unused-variable -Wno-unused-parameter -DTROPNLL2DP" ;
		:f90_compiler_version = "GNU Fortran (GCC) 4.8.5 20150623 (Red Hat 4.8.5-44)" ;
		:f90_compiler_flags = "-gdwarf-3 -O2 -fPIC -cpp -ffpe-trap=invalid -fno-range-check -frecursive -fimplicit-none -ffree-line-length-none -DTROPNLL2DP -Wuninitialized -Wtabs" ;
		:build_date = "2023-09-28T07:04:00Z" ;
		:revision_control_identifier = "d084fd110d84" ;
		:geolocation_grid_from_band = 4 ;
		:identifier_product_doi = "N/A" ;
		:identifier_product_doi_authority = "http://dx.doi.org/" ;
		:algorithm_version = "1.6.0" ;
		:title = "TROPOMI/S5P NO2 5-minute L2 Swath 5.5x3.5km" ;
		:processing_status = "NRTI-processing product" ;
		:product_version = "2.4.0" ;
		:Status_MET_2D = "Nominal" ;
		:Status_NISE__ = "Retired" ;
		:Status_CTMFCT = "Nominal" ;

group: PRODUCT {
  dimensions:
  	scanline = 372 ;
  	ground_pixel = 450 ;
  	corner = 4 ;
  	time = 1 ;
  	polynomial_exponents = 6 ;
  	intensity_offset_polynomial_exponents = 1 ;
  	layer = 34 ;
  	vertices = 2 ;
  variables:
  	int scanline(scanline) ;
  		scanline:units = "1" ;
  		scanline:axis = "Y" ;
  		scanline:long_name = "along-track dimension index" ;
  		scanline:comment = "This coordinate variable defines the indices along track; index starts at 0" ;
  		scanline:_FillValue = -2147483647 ;
  	int ground_pixel(ground_pixel) ;
  		ground_pixel:units = "1" ;
  		ground_pixel:axis = "X" ;
  		ground_pixel:long_name = "across-track dimension index" ;
  		ground_pixel:comment = "This coordinate variable defines the indices across track, from west to east; index starts at 0" ;
  		ground_pixel:_FillValue = -2147483647 ;
  	int time(time) ;
  		time:units = "seconds since 2010-01-01 00:00:00" ;
  		time:standard_name = "time" ;
  		time:axis = "T" ;
  		time:long_name = "reference time for the measurements" ;
  		time:comment = "The time in this variable corresponds to the time in the time_reference global attribute" ;
  		time:_FillValue = -2147483647 ;
  	int corner(corner) ;
  		corner:units = "1" ;
  		corner:long_name = "pixel corner index" ;
  		corner:comment = "This coordinate variable defines the indices for the pixel corners; index starts at 0 (counter-clockwise, starting from south-western corner of the pixel in ascending part of the orbit)" ;
  		corner:_FillValue = -2147483647 ;
  	int polynomial_exponents(polynomial_exponents) ;
  		polynomial_exponents:units = "1" ;
  		polynomial_exponents:long_name = "Polynomial exponents for background polynomial" ;
  		polynomial_exponents:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/polynomial_coefficients" ;
  		polynomial_exponents:_FillValue = -2147483647 ;
  	int intensity_offset_polynomial_exponents(intensity_offset_polynomial_exponents) ;
  		intensity_offset_polynomial_exponents:units = "1" ;
  		intensity_offset_polynomial_exponents:long_name = "Polynomial exponents for intensity offset" ;
  		intensity_offset_polynomial_exponents:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/polynomial_coefficients" ;
  		intensity_offset_polynomial_exponents:_FillValue = -2147483647 ;
  	int layer(layer) ;
  		layer:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
  		layer:units = "1" ;
  		layer:long_name = "TM5 atmospheric layer numbers" ;
  		layer:positive = "down" ;
  		layer:axis = "Z" ;
  		layer:formula_terms = "ap: tm5_constant_a b: tm5_constant_b ps: /PRODUCT/SUPPORT_DATA/INPUT_DATA/surface_pressure" ;
  		layer:comment = "p(t, k, j, i, l) = ap(k, l) + b(k, l)*ps(t, j, i); k from surface to top of atmosphere; l=0 for base of layer, l=1 for top of layer." ;
  		layer:_FillValue = -2147483647 ;
  	int vertices(vertices) ;
  		vertices:units = "1" ;
  		vertices:long_name = "TM5 atmospheric layer upper and lower bound indices" ;
  		vertices:_FillValue = -2147483647 ;
  	float latitude(time, scanline, ground_pixel) ;
  		latitude:long_name = "pixel center latitude" ;
  		latitude:units = "degrees_north" ;
  		latitude:standard_name = "latitude" ;
  		latitude:valid_min = -90.f ;
  		latitude:valid_max = 90.f ;
  		latitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/latitude_bounds" ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(time, scanline, ground_pixel) ;
  		longitude:long_name = "pixel center longitude" ;
  		longitude:units = "degrees_east" ;
  		longitude:standard_name = "longitude" ;
  		longitude:valid_min = -180.f ;
  		longitude:valid_max = 180.f ;
  		longitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/longitude_bounds" ;
  		longitude:_FillValue = 9.96921e+36f ;
  	int delta_time(time, scanline) ;
  		delta_time:long_name = "offset of start time of measurement relative to time_reference" ;
  		delta_time:units = "milliseconds since 2024-01-24 00:00:00" ;
  		delta_time:_FillValue = -2147483647 ;
  	string time_utc(time, scanline) ;
  		time_utc:long_name = "Time of observation as ISO 8601 date-time string" ;
  		string time_utc:_FillValue = "" ;
  	ubyte qa_value(time, scanline, ground_pixel) ;
  		qa_value:units = "1" ;
  		qa_value:scale_factor = 0.01f ;
  		qa_value:add_offset = 0.f ;
  		qa_value:valid_min = 0UB ;
  		qa_value:valid_max = 100UB ;
  		qa_value:long_name = "data quality value" ;
  		qa_value:comment = "A continuous quality descriptor, varying between 0 (no data) and 1 (full quality data). Recommend to ignore data with qa_value < 0.5" ;
  		qa_value:coordinates = "longitude latitude" ;
  		qa_value:_FillValue = 255UB ;
  	float nitrogendioxide_tropospheric_column(time, scanline, ground_pixel) ;
  		nitrogendioxide_tropospheric_column:units = "mol m-2" ;
  		nitrogendioxide_tropospheric_column:standard_name = "troposphere_mole_content_of_nitrogen_dioxide" ;
  		nitrogendioxide_tropospheric_column:long_name = "Tropospheric vertical column of nitrogen dioxide" ;
  		nitrogendioxide_tropospheric_column:coordinates = "longitude latitude" ;
  		nitrogendioxide_tropospheric_column:ancillary_variables = "nitrogendioxide_tropospheric_column_precision air_mass_factor_troposphere air_mass_factor_total averaging_kernel" ;
  		nitrogendioxide_tropospheric_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
  		nitrogendioxide_tropospheric_column:_FillValue = 9.96921e+36f ;
  	float nitrogendioxide_tropospheric_column_precision(time, scanline, ground_pixel) ;
  		nitrogendioxide_tropospheric_column_precision:units = "mol m-2" ;
  		nitrogendioxide_tropospheric_column_precision:standard_name = "troposphere_mole_content_of_nitrogen_dioxide standard_error" ;
  		nitrogendioxide_tropospheric_column_precision:long_name = "Precision of the tropospheric vertical column of nitrogen dioxide" ;
  		nitrogendioxide_tropospheric_column_precision:coordinates = "longitude latitude" ;
  		nitrogendioxide_tropospheric_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
  		nitrogendioxide_tropospheric_column_precision:_FillValue = 9.96921e+36f ;
  	float nitrogendioxide_tropospheric_column_precision_kernel(time, scanline, ground_pixel) ;
  		nitrogendioxide_tropospheric_column_precision_kernel:units = "mol m-2" ;
  		nitrogendioxide_tropospheric_column_precision_kernel:standard_name = "troposphere_mole_content_of_nitrogen_dioxide standard_error" ;
  		nitrogendioxide_tropospheric_column_precision_kernel:long_name = "Precision of the tropospheric vertical column of nitrogen dioxide when applying the averaging kernel" ;
  		nitrogendioxide_tropospheric_column_precision_kernel:coordinates = "longitude latitude" ;
  		nitrogendioxide_tropospheric_column_precision_kernel:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
  		nitrogendioxide_tropospheric_column_precision_kernel:_FillValue = 9.96921e+36f ;
  	float averaging_kernel(time, scanline, ground_pixel, layer) ;
  		averaging_kernel:units = "1" ;
  		averaging_kernel:long_name = "Averaging kernel" ;
  		averaging_kernel:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  		averaging_kernel:ancillary_variables = "tm5_constant_a tm5_constant_b tm5_tropopause_layer_index /PRODUCT/SUPPORT_DATA/INPUT_DATA/surface_pressure" ;
  		averaging_kernel:_FillValue = 9.96921e+36f ;
  	float air_mass_factor_troposphere(time, scanline, ground_pixel) ;
  		air_mass_factor_troposphere:units = "1" ;
  		air_mass_factor_troposphere:long_name = "Tropospheric air mass factor" ;
  		air_mass_factor_troposphere:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  		air_mass_factor_troposphere:ancillary_variables = "tm5_tropopause_layer_index" ;
  		air_mass_factor_troposphere:_FillValue = 9.96921e+36f ;
  	float air_mass_factor_total(time, scanline, ground_pixel) ;
  		air_mass_factor_total:units = "1" ;
  		air_mass_factor_total:long_name = "Total air mass factor" ;
  		air_mass_factor_total:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  		air_mass_factor_total:_FillValue = 9.96921e+36f ;
  	int tm5_tropopause_layer_index(time, scanline, ground_pixel) ;
  		tm5_tropopause_layer_index:units = "1" ;
  		tm5_tropopause_layer_index:long_name = "TM5 layer index of the highest layer in the tropopause" ;
  		tm5_tropopause_layer_index:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  		tm5_tropopause_layer_index:ancillary_variables = "tm5_constant_a tm5_constant_b /PRODUCT/SUPPORT_DATA/INPUT_DATA/surface_pressure" ;
  		tm5_tropopause_layer_index:_FillValue = -2147483647 ;
  	float tm5_constant_a(layer, vertices) ;
  		tm5_constant_a:units = "Pa" ;
  		tm5_constant_a:long_name = "TM5 hybrid A coefficient at upper and lower interface levels" ;
  		tm5_constant_a:_FillValue = 9.96921e+36f ;
  	float tm5_constant_b(layer, vertices) ;
  		tm5_constant_b:units = "1" ;
  		tm5_constant_b:long_name = "TM5 hybrid B coefficient at upper and lower interface levels" ;
  		tm5_constant_b:_FillValue = 9.96921e+36f ;

  group: SUPPORT_DATA {

    group: GEOLOCATIONS {
      variables:
      	float satellite_latitude(time, scanline) ;
      		satellite_latitude:long_name = "sub satellite latitude" ;
      		satellite_latitude:units = "degrees_north" ;
      		satellite_latitude:comment = "Latitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_latitude:valid_min = -90.f ;
      		satellite_latitude:valid_max = 90.f ;
      		satellite_latitude:_FillValue = 9.96921e+36f ;
      	float satellite_longitude(time, scanline) ;
      		satellite_longitude:long_name = "satellite_longitude" ;
      		satellite_longitude:units = "degrees_east" ;
      		satellite_longitude:comment = "Longitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_longitude:valid_min = -180.f ;
      		satellite_longitude:valid_max = 180.f ;
      		satellite_longitude:_FillValue = 9.96921e+36f ;
      	float satellite_altitude(time, scanline) ;
      		satellite_altitude:long_name = "satellite altitude" ;
      		satellite_altitude:units = "m" ;
      		satellite_altitude:comment = "The altitude of the satellite with respect to the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_altitude:valid_min = 700000.f ;
      		satellite_altitude:valid_max = 900000.f ;
      		satellite_altitude:_FillValue = 9.96921e+36f ;
      	float satellite_orbit_phase(time, scanline) ;
      		satellite_orbit_phase:long_name = "fractional satellite orbit phase" ;
      		satellite_orbit_phase:units = "1" ;
      		satellite_orbit_phase:comment = "Relative offset [0.0, ..., 1.0] of the measurement in the orbit" ;
      		satellite_orbit_phase:valid_min = -0.02f ;
      		satellite_orbit_phase:valid_max = 1.02f ;
      		satellite_orbit_phase:_FillValue = 9.96921e+36f ;
      	float solar_zenith_angle(time, scanline, ground_pixel) ;
      		solar_zenith_angle:long_name = "solar zenith angle" ;
      		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
      		solar_zenith_angle:units = "degree" ;
      		solar_zenith_angle:valid_min = 0.f ;
      		solar_zenith_angle:valid_max = 180.f ;
      		solar_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_zenith_angle:comment = "Solar zenith angle at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      		solar_zenith_angle:_FillValue = 9.96921e+36f ;
      	float solar_azimuth_angle(time, scanline, ground_pixel) ;
      		solar_azimuth_angle:long_name = "solar azimuth angle" ;
      		solar_azimuth_angle:standard_name = "solar_azimuth_angle" ;
      		solar_azimuth_angle:units = "degree" ;
      		solar_azimuth_angle:valid_min = -180.f ;
      		solar_azimuth_angle:valid_max = 180.f ;
      		solar_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_azimuth_angle:comment = "Solar azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = +/-180, West = -90)" ;
      		solar_azimuth_angle:_FillValue = 9.96921e+36f ;
      	float viewing_zenith_angle(time, scanline, ground_pixel) ;
      		viewing_zenith_angle:long_name = "viewing zenith angle" ;
      		viewing_zenith_angle:standard_name = "viewing_zenith_angle" ;
      		viewing_zenith_angle:units = "degree" ;
      		viewing_zenith_angle:valid_min = 0.f ;
      		viewing_zenith_angle:valid_max = 180.f ;
      		viewing_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_zenith_angle:comment = "Zenith angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      		viewing_zenith_angle:_FillValue = 9.96921e+36f ;
      	float viewing_azimuth_angle(time, scanline, ground_pixel) ;
      		viewing_azimuth_angle:long_name = "viewing azimuth angle" ;
      		viewing_azimuth_angle:standard_name = "viewing_azimuth_angle" ;
      		viewing_azimuth_angle:units = "degree" ;
      		viewing_azimuth_angle:valid_min = -180.f ;
      		viewing_azimuth_angle:valid_max = 180.f ;
      		viewing_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_azimuth_angle:comment = "Satellite azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = +/-180, West = -90)" ;
      		viewing_azimuth_angle:_FillValue = 9.96921e+36f ;
      	float latitude_bounds(time, scanline, ground_pixel, corner) ;
      		latitude_bounds:_FillValue = 9.96921e+36f ;
      	float longitude_bounds(time, scanline, ground_pixel, corner) ;
      		longitude_bounds:_FillValue = 9.96921e+36f ;
      	ubyte geolocation_flags(time, scanline, ground_pixel) ;
      		geolocation_flags:_FillValue = 255UB ;
      		geolocation_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		geolocation_flags:flag_masks = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 128UB ;
      		geolocation_flags:flag_meanings = "no_error solar_eclipse sun_glint_possible descending night geo_boundary_crossing spacecraft_manoeuvre geolocation_error" ;
      		geolocation_flags:flag_values = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 128UB ;
      		geolocation_flags:long_name = "geolocation flags" ;
      		geolocation_flags:max_val = 254UB ;
      		geolocation_flags:min_val = 0UB ;
      		geolocation_flags:units = "1" ;
      } // group GEOLOCATIONS

    group: DETAILED_RESULTS {
      variables:
      	uint processing_quality_flags(time, scanline, ground_pixel) ;
      		processing_quality_flags:long_name = "Processing quality flags" ;
      		processing_quality_flags:comment = "Flags indicating conditions that affect quality of the retrieval." ;
      		processing_quality_flags:flag_meanings = "success radiance_missing irradiance_missing input_spectrum_missing reflectance_range_error ler_range_error snr_range_error sza_range_error vza_range_error lut_range_error ozone_range_error wavelength_offset_error initialization_error memory_error assertion_error io_error numerical_error lut_error ISRF_error convergence_error cloud_filter_convergence_error max_iteration_convergence_error aot_lower_boundary_convergence_error other_boundary_convergence_error geolocation_error ch4_noscat_zero_error h2o_noscat_zero_error max_optical_thickness_error aerosol_boundary_error boundary_hit_error chi2_error svd_error dfs_error radiative_transfer_error optimal_estimation_error profile_error cloud_error model_error number_of_input_data_points_too_low_error cloud_pressure_spread_too_low_error cloud_too_low_level_error generic_range_error generic_exception input_spectrum_alignment_error abort_error wrong_input_type_error wavelength_calibration_error coregistration_error slant_column_density_error airmass_factor_error vertical_column_density_error signal_to_noise_ratio_error configuration_error key_error saturation_error max_num_outlier_exceeded_error solar_eclipse_filter cloud_filter altitude_consistency_filter altitude_roughness_filter sun_glint_filter mixed_surface_type_filter snow_ice_filter aai_filter cloud_fraction_fresco_filter aai_scene_albedo_filter small_pixel_radiance_std_filter cloud_fraction_viirs_filter cirrus_reflectance_viirs_filter cf_viirs_swir_ifov_filter cf_viirs_swir_ofova_filter cf_viirs_swir_ofovb_filter cf_viirs_swir_ofovc_filter cf_viirs_nir_ifov_filter cf_viirs_nir_ofova_filter cf_viirs_nir_ofovb_filter cf_viirs_nir_ofovc_filter refl_cirrus_viirs_swir_filter refl_cirrus_viirs_nir_filter diff_refl_cirrus_viirs_filter ch4_noscat_ratio_filter ch4_noscat_ratio_std_filter h2o_noscat_ratio_filter h2o_noscat_ratio_std_filter diff_psurf_fresco_ecmwf_filter psurf_fresco_stdv_filter ocean_filter time_range_filter pixel_or_scanline_index_filter geographic_region_filter internal_cloud_mask_filter input_spectrum_warning wavelength_calibration_warning extrapolation_warning sun_glint_warning south_atlantic_anomaly_warning sun_glint_correction snow_ice_warning cloud_warning AAI_warning pixel_level_input_data_missing data_range_warning low_cloud_fraction_warning altitude_consistency_warning signal_to_noise_ratio_warning deconvolution_warning so2_volcanic_origin_likely_warning so2_volcanic_origin_certain_warning interpolation_warning saturation_warning high_sza_warning cloud_retrieval_warning cloud_inhomogeneity_warning thermal_instability_warning" ;
      		processing_quality_flags:flag_masks = 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U, 67108864U, 134217728U, 268435456U, 536870912U, 1073741824U ;
      		processing_quality_flags:flag_values = 0U, 1U, 2U, 3U, 4U, 5U, 6U, 7U, 8U, 9U, 10U, 11U, 12U, 13U, 14U, 15U, 16U, 17U, 18U, 19U, 20U, 21U, 22U, 23U, 24U, 25U, 26U, 27U, 28U, 29U, 30U, 31U, 32U, 33U, 34U, 35U, 36U, 37U, 38U, 39U, 40U, 41U, 42U, 43U, 44U, 45U, 46U, 47U, 48U, 49U, 50U, 51U, 52U, 53U, 54U, 55U, 64U, 65U, 66U, 67U, 68U, 69U, 70U, 71U, 72U, 73U, 74U, 75U, 76U, 77U, 78U, 79U, 80U, 81U, 82U, 83U, 84U, 85U, 86U, 87U, 88U, 89U, 90U, 91U, 92U, 93U, 94U, 95U, 96U, 97U, 98U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U, 67108864U, 134217728U, 268435456U, 536870912U, 1073741824U ;
      		processing_quality_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		processing_quality_flags:_FillValue = 4294967295U ;
      	ushort number_of_spectral_points_in_retrieval(time, scanline, ground_pixel) ;
      		number_of_spectral_points_in_retrieval:long_name = "Number of spectral points used in the retrieval" ;
      		number_of_spectral_points_in_retrieval:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		number_of_spectral_points_in_retrieval:_FillValue = 65535US ;
      	int number_of_iterations(time, scanline, ground_pixel) ;
      		number_of_iterations:long_name = "number of iterations" ;
      		number_of_iterations:units = "1" ;
      		number_of_iterations:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		number_of_iterations:_FillValue = -2147483647 ;
      	float wavelength_calibration_offset(time, scanline, ground_pixel) ;
      		wavelength_calibration_offset:long_name = "radiance wavelength offset" ;
      		wavelength_calibration_offset:units = "nm" ;
      		wavelength_calibration_offset:wavelength_fit_window_start = 405. ;
      		wavelength_calibration_offset:wavelength_fit_window_end = 465. ;
      		wavelength_calibration_offset:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_offset:ancillary_variables = "wavelength_calibration_offset_precision" ;
      		wavelength_calibration_offset:comment = "True wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
      		wavelength_calibration_offset:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_offset_precision(time, scanline, ground_pixel) ;
      		wavelength_calibration_offset_precision:long_name = "radiance wavelength offset precision" ;
      		wavelength_calibration_offset_precision:units = "nm" ;
      		wavelength_calibration_offset_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_offset_precision:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_stretch(time, scanline, ground_pixel) ;
      		wavelength_calibration_stretch:long_name = "radiance wavelength stretch" ;
      		wavelength_calibration_stretch:units = "1" ;
      		wavelength_calibration_stretch:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_stretch:ancillary_variables = "wavelength_calibration_stretch_precision" ;
      		wavelength_calibration_stretch:comment = "True wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
      		wavelength_calibration_stretch:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_stretch_precision(time, scanline, ground_pixel) ;
      		wavelength_calibration_stretch_precision:long_name = "radiance wavelength stretch precision" ;
      		wavelength_calibration_stretch_precision:units = "1" ;
      		wavelength_calibration_stretch_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_stretch_precision:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_chi_square(time, scanline, ground_pixel) ;
      		wavelength_calibration_chi_square:long_name = "radiance wavelength calibration chi square" ;
      		wavelength_calibration_chi_square:units = "1" ;
      		wavelength_calibration_chi_square:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_chi_square:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_irradiance_offset(time, ground_pixel) ;
      		wavelength_calibration_irradiance_offset:long_name = "irradiance wavelength offset" ;
      		wavelength_calibration_irradiance_offset:units = "nm" ;
      		wavelength_calibration_irradiance_offset:wavelength_fit_window_start = 405. ;
      		wavelength_calibration_irradiance_offset:wavelength_fit_window_end = 465. ;
      		wavelength_calibration_irradiance_offset:ancillary_variables = "wavelength_calibration_irradiance_offset_precision" ;
      		wavelength_calibration_irradiance_offset:comment = "True wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
      		wavelength_calibration_irradiance_offset:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_irradiance_offset_precision(time, ground_pixel) ;
      		wavelength_calibration_irradiance_offset_precision:long_name = "irradiance wavelength offset precision" ;
      		wavelength_calibration_irradiance_offset_precision:units = "nm" ;
      		wavelength_calibration_irradiance_offset_precision:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_irradiance_chi_square(time, ground_pixel) ;
      		wavelength_calibration_irradiance_chi_square:long_name = "irradiance wavelength calibration chi squared" ;
      		wavelength_calibration_irradiance_chi_square:units = "1" ;
      		wavelength_calibration_irradiance_chi_square:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_stratospheric_column(time, scanline, ground_pixel) ;
      		nitrogendioxide_stratospheric_column:units = "mol m-2" ;
      		nitrogendioxide_stratospheric_column:standard_name = "stratosphere_mole_content_of_nitrogen_dioxide" ;
      		nitrogendioxide_stratospheric_column:long_name = "Stratospheric vertical column of nitrogen dioxide, derived from the TM5-MP vertical profiles" ;
      		nitrogendioxide_stratospheric_column:coordinates = "longitude latitude" ;
      		nitrogendioxide_stratospheric_column:ancillary_variables = "nitrogendioxide_stratospheric_column_precision air_mass_factor_stratosphere /PRODUCT/air_mass_factor_total /PRODUCT/averaging_kernel" ;
      		nitrogendioxide_stratospheric_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_stratospheric_column:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_stratospheric_column_precision(time, scanline, ground_pixel) ;
      		nitrogendioxide_stratospheric_column_precision:units = "mol m-2" ;
      		nitrogendioxide_stratospheric_column_precision:standard_name = "stratosphere_mole_content_of_nitrogen_dioxide standard_error" ;
      		nitrogendioxide_stratospheric_column_precision:long_name = "Precision of stratospheric vertical column of nitrogen dioxide" ;
      		nitrogendioxide_stratospheric_column_precision:coordinates = "longitude latitude" ;
      		nitrogendioxide_stratospheric_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_stratospheric_column_precision:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_total_column(time, scanline, ground_pixel) ;
      		nitrogendioxide_total_column:units = "mol m-2" ;
      		nitrogendioxide_total_column:proposed_standard_name = "atmosphere_mole_content_of_nitrogen_dioxide" ;
      		nitrogendioxide_total_column:long_name = "Total vertical column of nitrogen dioxide derived from the total slant column and TM5 profile in stratosphere and troposphere" ;
      		nitrogendioxide_total_column:coordinates = "longitude latitude" ;
      		nitrogendioxide_total_column:ancillary_variables = "nitrogendioxide_total_column_precision /PRODUCT/averaging_kernel" ;
      		nitrogendioxide_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_total_column:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_total_column_precision(time, scanline, ground_pixel) ;
      		nitrogendioxide_total_column_precision:units = "mol m-2" ;
      		nitrogendioxide_total_column_precision:proposed_standard_name = "atmosphere_mole_content_of_nitrogen_dioxide standard_error" ;
      		nitrogendioxide_total_column_precision:long_name = "Precision of the total vertical column of nitrogen dioxide derived from the total slant column and TM5 profile in stratosphere and troposphere" ;
      		nitrogendioxide_total_column_precision:coordinates = "longitude latitude" ;
      		nitrogendioxide_total_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_total_column_precision:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_total_column_precision_kernel(time, scanline, ground_pixel) ;
      		nitrogendioxide_total_column_precision_kernel:units = "mol m-2" ;
      		nitrogendioxide_total_column_precision_kernel:proposed_standard_name = "atmosphere_mole_content_of_nitrogen_dioxide standard_error" ;
      		nitrogendioxide_total_column_precision_kernel:long_name = "Precision of the total vertical column of nitrogen dioxide derived from the total slant column and TM5 profile in stratosphere and troposphere, when the averaging kernel is applied" ;
      		nitrogendioxide_total_column_precision_kernel:coordinates = "longitude latitude" ;
      		nitrogendioxide_total_column_precision_kernel:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_total_column_precision_kernel:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_summed_total_column(time, scanline, ground_pixel) ;
      		nitrogendioxide_summed_total_column:units = "mol m-2" ;
      		nitrogendioxide_summed_total_column:proposed_standard_name = "atmosphere_mole_content_of_nitrogen_dioxide" ;
      		nitrogendioxide_summed_total_column:long_name = "Sum of the tropospheric and stratospheric vertical columns" ;
      		nitrogendioxide_summed_total_column:coordinates = "longitude latitude" ;
      		nitrogendioxide_summed_total_column:ancillary_variables = "nitrogendioxide_summed_total_column_precision" ;
      		nitrogendioxide_summed_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_summed_total_column:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_summed_total_column_precision(time, scanline, ground_pixel) ;
      		nitrogendioxide_summed_total_column_precision:units = "mol m-2" ;
      		nitrogendioxide_summed_total_column_precision:proposed_standard_name = "atmosphere_mole_content_of_nitrogen_dioxide standard_error" ;
      		nitrogendioxide_summed_total_column_precision:long_name = "Precision of the sum of the tropospheric and stratospheric vertical columns" ;
      		nitrogendioxide_summed_total_column_precision:coordinates = "longitude latitude" ;
      		nitrogendioxide_summed_total_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_summed_total_column_precision:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_slant_column_density(time, scanline, ground_pixel) ;
      		nitrogendioxide_slant_column_density:units = "mol m-2" ;
      		nitrogendioxide_slant_column_density:long_name = "NO2 slant column density" ;
      		nitrogendioxide_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		nitrogendioxide_slant_column_density:ancillary_variables = "nitrogendioxide_slant_column_density_precision" ;
      		nitrogendioxide_slant_column_density:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_slant_column_density:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_slant_column_density_precision(time, scanline, ground_pixel) ;
      		nitrogendioxide_slant_column_density_precision:units = "mol m-2" ;
      		nitrogendioxide_slant_column_density_precision:long_name = "NO2 slant column density precision" ;
      		nitrogendioxide_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		nitrogendioxide_slant_column_density_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_slant_column_density_precision:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_slant_column_density_stripe_amplitude(time, ground_pixel) ;
      		nitrogendioxide_slant_column_density_stripe_amplitude:units = "mol m-2" ;
      		nitrogendioxide_slant_column_density_stripe_amplitude:long_name = "Across-track NO2 slant column stripe offset, 7-day mean, determined over the Pacific Ocean" ;
      		nitrogendioxide_slant_column_density_stripe_amplitude:comment = "The stripe amplitude is subtracted from the NO2 slant column before the vertical columns are computed" ;
      		nitrogendioxide_slant_column_density_stripe_amplitude:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_slant_column_density_stripe_amplitude:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_geometric_column(time, scanline, ground_pixel) ;
      		nitrogendioxide_geometric_column:long_name = "Geometric vertical column geometric column of nitrogen dioxide" ;
      		nitrogendioxide_geometric_column:comment = "The geometric column (GCD) is the slant column (SCD) divided by geometric air-mass factor (AMFgeo)" ;
      		nitrogendioxide_geometric_column:units = "mol m-2" ;
      		nitrogendioxide_geometric_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_geometric_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		nitrogendioxide_geometric_column:ancillary_variables = "nitrogendioxide_geometric_column_precision" ;
      		nitrogendioxide_geometric_column:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_geometric_column_precision(time, scanline, ground_pixel) ;
      		nitrogendioxide_geometric_column_precision:long_name = "Precision of the geometric vertical column geometric column of nitrogen dioxide" ;
      		nitrogendioxide_geometric_column_precision:units = "mol m-2" ;
      		nitrogendioxide_geometric_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_geometric_column_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		nitrogendioxide_geometric_column_precision:_FillValue = 9.96921e+36f ;
      	float ozone_slant_column_density(time, scanline, ground_pixel) ;
      		ozone_slant_column_density:units = "mol m-2" ;
      		ozone_slant_column_density:long_name = "O3 slant column density" ;
      		ozone_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		ozone_slant_column_density:ancillary_variables = "ozone_slant_column_density_precision" ;
      		ozone_slant_column_density:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		ozone_slant_column_density:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		ozone_slant_column_density:_FillValue = 9.96921e+36f ;
      	float ozone_slant_column_density_precision(time, scanline, ground_pixel) ;
      		ozone_slant_column_density_precision:units = "mol m-2" ;
      		ozone_slant_column_density_precision:long_name = "O3 slant column density precision" ;
      		ozone_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		ozone_slant_column_density_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		ozone_slant_column_density_precision:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		ozone_slant_column_density_precision:_FillValue = 9.96921e+36f ;
      	float oxygen_oxygen_dimer_slant_column_density(time, scanline, ground_pixel) ;
      		oxygen_oxygen_dimer_slant_column_density:units = "mol2 m-5" ;
      		oxygen_oxygen_dimer_slant_column_density:long_name = "Slant column density of oxygen collision induced absorption" ;
      		oxygen_oxygen_dimer_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		oxygen_oxygen_dimer_slant_column_density:ancillary_variables = "oxygen_oxygen_dimer_slant_column_density_precision" ;
      		oxygen_oxygen_dimer_slant_column_density:multiplication_factor_to_convert_to_molecules2_percm5 = 3.62662e+37 ;
      		oxygen_oxygen_dimer_slant_column_density:_FillValue = 9.96921e+36f ;
      	float oxygen_oxygen_dimer_slant_column_density_precision(time, scanline, ground_pixel) ;
      		oxygen_oxygen_dimer_slant_column_density_precision:units = "mol2 m-5" ;
      		oxygen_oxygen_dimer_slant_column_density_precision:long_name = "Precision of the slant column density of oxygen collision induced absorption" ;
      		oxygen_oxygen_dimer_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		oxygen_oxygen_dimer_slant_column_density_precision:multiplication_factor_to_convert_to_molecules2_percm5 = 3.62662e+37 ;
      		oxygen_oxygen_dimer_slant_column_density_precision:_FillValue = 9.96921e+36f ;
      	float water_slant_column_density(time, scanline, ground_pixel) ;
      		water_slant_column_density:units = "mol m-2" ;
      		water_slant_column_density:long_name = "Water vapor slant column density" ;
      		water_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_slant_column_density:ancillary_variables = "water_slant_column_density_precision" ;
      		water_slant_column_density:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		water_slant_column_density:_FillValue = 9.96921e+36f ;
      	float water_slant_column_density_precision(time, scanline, ground_pixel) ;
      		water_slant_column_density_precision:units = "mol m-2" ;
      		water_slant_column_density_precision:long_name = "Precision of water vapor slant column density" ;
      		water_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_slant_column_density_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		water_slant_column_density_precision:_FillValue = 9.96921e+36f ;
      	float water_liquid_slant_column_density(time, scanline, ground_pixel) ;
      		water_liquid_slant_column_density:units = "m" ;
      		water_liquid_slant_column_density:long_name = "Liquid water column" ;
      		water_liquid_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_liquid_slant_column_density:ancillary_variables = "water_liquid_slant_column_density_precision" ;
      		water_liquid_slant_column_density:_FillValue = 9.96921e+36f ;
      	float water_liquid_slant_column_density_precision(time, scanline, ground_pixel) ;
      		water_liquid_slant_column_density_precision:units = "m" ;
      		water_liquid_slant_column_density_precision:long_name = "Precision of liquid water column" ;
      		water_liquid_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_liquid_slant_column_density_precision:_FillValue = 9.96921e+36f ;
      	float ring_coefficient(time, scanline, ground_pixel) ;
      		ring_coefficient:units = "1" ;
      		ring_coefficient:long_name = "Fit coefficient of the Ring effect" ;
      		ring_coefficient:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		ring_coefficient:ancillary_variables = "ring_coefficient_precision" ;
      		ring_coefficient:_FillValue = 9.96921e+36f ;
      	float ring_coefficient_precision(time, scanline, ground_pixel) ;
      		ring_coefficient_precision:units = "1" ;
      		ring_coefficient_precision:long_name = "Precision of fit coefficient of the Ring effect" ;
      		ring_coefficient_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		ring_coefficient_precision:_FillValue = 9.96921e+36f ;
      	float polynomial_coefficients(time, scanline, ground_pixel, polynomial_exponents) ;
      		polynomial_coefficients:units = "1" ;
      		polynomial_coefficients:long_name = "Polynomial coefficients of the DOAS fit" ;
      		polynomial_coefficients:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		polynomial_coefficients:ancillary_variables = "polynomial_coefficients_precision" ;
      		polynomial_coefficients:_FillValue = 9.96921e+36f ;
      	float polynomial_coefficients_precision(time, scanline, ground_pixel, polynomial_exponents) ;
      		polynomial_coefficients_precision:units = "1" ;
      		polynomial_coefficients_precision:long_name = "Precision of the polynomial coefficients of the DOAS fit" ;
      		polynomial_coefficients_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		polynomial_coefficients_precision:_FillValue = 9.96921e+36f ;
      	float intensity_offset_coefficients(time, scanline, ground_pixel, intensity_offset_polynomial_exponents) ;
      		intensity_offset_coefficients:units = "1" ;
      		intensity_offset_coefficients:long_name = "Polynomial coefficients of the intensity offset" ;
      		intensity_offset_coefficients:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		intensity_offset_coefficients:ancillary_variables = "polynomial_coefficients_precision" ;
      		intensity_offset_coefficients:_FillValue = 9.96921e+36f ;
      	float intensity_offset_coefficients_precision(time, scanline, ground_pixel, intensity_offset_polynomial_exponents) ;
      		intensity_offset_coefficients_precision:units = "1" ;
      		intensity_offset_coefficients_precision:long_name = "Precision of the polynomial coefficients of the intensity offset" ;
      		intensity_offset_coefficients_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		intensity_offset_coefficients_precision:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_crb_nitrogendioxide_window(time, scanline, ground_pixel) ;
      		cloud_fraction_crb_nitrogendioxide_window:proposed_standard_name = "effective_cloud_area_fraction_assuming_fixed_cloud_albedo" ;
      		cloud_fraction_crb_nitrogendioxide_window:units = "1" ;
      		cloud_fraction_crb_nitrogendioxide_window:long_name = "Cloud fraction at 440 nm for NO2 retrieval" ;
      		cloud_fraction_crb_nitrogendioxide_window:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_crb_nitrogendioxide_window:radiation_wavelength = 440.f ;
      		cloud_fraction_crb_nitrogendioxide_window:assumed_cloud_albedo = 0.8f ;
      		cloud_fraction_crb_nitrogendioxide_window:ancillary_variables = "cloud_radiance_fraction_nitrogendioxide_window /PRODUCT/SUPPORT_DATA/INPUT_DATA/cloud_pressure_crb" ;
      		cloud_fraction_crb_nitrogendioxide_window:_FillValue = 9.96921e+36f ;
      	float cloud_radiance_fraction_nitrogendioxide_window(time, scanline, ground_pixel) ;
      		cloud_radiance_fraction_nitrogendioxide_window:units = "1" ;
      		cloud_radiance_fraction_nitrogendioxide_window:long_name = "Cloud radiance fraction at 440 nm for NO2 retrieval" ;
      		cloud_radiance_fraction_nitrogendioxide_window:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_radiance_fraction_nitrogendioxide_window:radiation_wavelength = 440.f ;
      		cloud_radiance_fraction_nitrogendioxide_window:assumed_cloud_albedo = 0.8f ;
      		cloud_radiance_fraction_nitrogendioxide_window:ancillary_variables = "cloud_fraction_crb_nitrogendioxide_window /PRODUCT/SUPPORT_DATA/INPUT_DATA/cloud_pressure_crb" ;
      		cloud_radiance_fraction_nitrogendioxide_window:_FillValue = 9.96921e+36f ;
      	float chi_square(time, scanline, ground_pixel) ;
      		chi_square:units = "1" ;
      		chi_square:long_name = "Chi squared of fit" ;
      		chi_square:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		chi_square:ancillary_variables = "number_of_spectral_points_in_retrieval degrees_of_freedom" ;
      		chi_square:_FillValue = 9.96921e+36f ;
      	float root_mean_square_error_of_fit(time, scanline, ground_pixel) ;
      		root_mean_square_error_of_fit:units = "1" ;
      		root_mean_square_error_of_fit:long_name = "Root mean square residual of the fit" ;
      		root_mean_square_error_of_fit:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		root_mean_square_error_of_fit:ancillary_variables = "number_of_spectral_points_in_retrieval" ;
      		root_mean_square_error_of_fit:_FillValue = 9.96921e+36f ;
      	float degrees_of_freedom(time, scanline, ground_pixel) ;
      		degrees_of_freedom:units = "1" ;
      		degrees_of_freedom:long_name = "Degrees of freedom from slant column fit" ;
      		degrees_of_freedom:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		degrees_of_freedom:ancillary_variables = "number_of_spectral_points_in_retrieval" ;
      		degrees_of_freedom:_FillValue = 9.96921e+36f ;
      	float air_mass_factor_stratosphere(time, scanline, ground_pixel) ;
      		air_mass_factor_stratosphere:units = "1" ;
      		air_mass_factor_stratosphere:long_name = "Stratospheric air mass factor" ;
      		air_mass_factor_stratosphere:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		air_mass_factor_stratosphere:ancillary_variables = "/PRODUCT/tm5_tropopause_layer_index" ;
      		air_mass_factor_stratosphere:_FillValue = 9.96921e+36f ;
      	float air_mass_factor_cloudy(time, scanline, ground_pixel) ;
      		air_mass_factor_cloudy:units = "1" ;
      		air_mass_factor_cloudy:long_name = "Air mass factor for the cloud-covered part of the scene" ;
      		air_mass_factor_cloudy:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		air_mass_factor_cloudy:ancillary_variables = "tm5_tropopause_layer_index" ;
      		air_mass_factor_cloudy:_FillValue = 9.96921e+36f ;
      	float air_mass_factor_clear(time, scanline, ground_pixel) ;
      		air_mass_factor_clear:units = "1" ;
      		air_mass_factor_clear:long_name = "Air mass factor for the cloud-free part of the scene" ;
      		air_mass_factor_clear:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		air_mass_factor_clear:ancillary_variables = "tm5_tropopause_layer_index" ;
      		air_mass_factor_clear:_FillValue = 9.96921e+36f ;
      	float nitrogendioxide_ghost_column(time, scanline, ground_pixel) ;
      		nitrogendioxide_ghost_column:units = "mol m-2" ;
      		nitrogendioxide_ghost_column:long_name = "Ghost column NO2: modelled NO2 column below the cloud top" ;
      		nitrogendioxide_ghost_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		nitrogendioxide_ghost_column:ancillary_variables = "/PRODUCT/SUPPORT_DATA/INPUT_DATA/cloud_pressure_crb" ;
      		nitrogendioxide_ghost_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      		nitrogendioxide_ghost_column:_FillValue = 9.96921e+36f ;
      	ubyte cloud_selection_flag(time, scanline, ground_pixel) ;
      		cloud_selection_flag:units = "1" ;
      		cloud_selection_flag:long_name = "Cloud product selection flag" ;
      		cloud_selection_flag:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_selection_flag:flag_values = 0UB, 1UB, 2UB, 4UB, 8UB ;
      		cloud_selection_flag:flag_meanings = "None FRESCO O22CLD CLOUD_ forced_selection" ;
      		cloud_selection_flag:flag_masks = 7UB, 7UB, 7UB, 7UB, 8UB ;
      		cloud_selection_flag:_FillValue = 255UB ;

      group: O22CLD {
        variables:
        	float o22cld_cloud_fraction_crb(time, scanline, ground_pixel) ;
        		o22cld_cloud_fraction_crb:units = "1" ;
        		o22cld_cloud_fraction_crb:long_name = "effective_cloud_area_fraction_assuming_fixed_cloud_albedo" ;
        		o22cld_cloud_fraction_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_fraction_crb:ancillary_variables = "o22cld_cloud_fraction_crb_precision" ;
        		o22cld_cloud_fraction_crb:_FillValue = 9.96921e+36f ;
        	float o22cld_cloud_fraction_crb_precision(time, scanline, ground_pixel) ;
        		o22cld_cloud_fraction_crb_precision:units = "1" ;
        		o22cld_cloud_fraction_crb_precision:long_name = "effective_cloud_area_fraction_assuming_fixed_cloud_albedo standard_error" ;
        		o22cld_cloud_fraction_crb_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_fraction_crb_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_cloud_pressure_crb(time, scanline, ground_pixel) ;
        		o22cld_cloud_pressure_crb:units = "Pa" ;
        		o22cld_cloud_pressure_crb:long_name = "air_pressure_at_cloud_optical_centroid" ;
        		o22cld_cloud_pressure_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_pressure_crb:ancillary_variables = "o22cld_cloud_pressure_crb_precision" ;
        		o22cld_cloud_pressure_crb:_FillValue = 9.96921e+36f ;
        	float o22cld_cloud_pressure_crb_precision(time, scanline, ground_pixel) ;
        		o22cld_cloud_pressure_crb_precision:units = "Pa" ;
        		o22cld_cloud_pressure_crb_precision:long_name = "air_pressure_at_cloud_optical_centroid standard_error" ;
        		o22cld_cloud_pressure_crb_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_pressure_crb_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_cloud_height_crb(time, scanline, ground_pixel) ;
        		o22cld_cloud_height_crb:units = "m" ;
        		o22cld_cloud_height_crb:long_name = "height_of_cloud_optical_centroid" ;
        		o22cld_cloud_height_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_height_crb:ancillary_variables = "o22cld_cloud_height_crb_precision" ;
        		o22cld_cloud_height_crb:_FillValue = 9.96921e+36f ;
        	float o22cld_cloud_height_crb_precision(time, scanline, ground_pixel) ;
        		o22cld_cloud_height_crb_precision:units = "m" ;
        		o22cld_cloud_height_crb_precision:long_name = "height_of_cloud_optical_centroid standard_error" ;
        		o22cld_cloud_height_crb_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_height_crb_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_cloud_albedo_crb(time, scanline, ground_pixel) ;
        		o22cld_cloud_albedo_crb:units = "1" ;
        		o22cld_cloud_albedo_crb:standard_name = "cloud_albedo" ;
        		o22cld_cloud_albedo_crb:long_name = "cloud albedo" ;
        		o22cld_cloud_albedo_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_cloud_albedo_crb:_FillValue = 9.96921e+36f ;
        	float o22cld_scene_albedo(time, scanline, ground_pixel) ;
        		o22cld_scene_albedo:units = "1" ;
        		o22cld_scene_albedo:long_name = "cloud_albedo_assuming_completely_cloudy_sky" ;
        		o22cld_scene_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_scene_albedo:ancillary_variables = "o22cld_scene_albedo_precision" ;
        		o22cld_scene_albedo:_FillValue = 9.96921e+36f ;
        	float o22cld_scene_albedo_precision(time, scanline, ground_pixel) ;
        		o22cld_scene_albedo_precision:units = "1" ;
        		o22cld_scene_albedo_precision:long_name = "cloud_albedo_assuming_completely_cloudy_sky standard_error" ;
        		o22cld_scene_albedo_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_scene_albedo_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_apparent_scene_pressure(time, scanline, ground_pixel) ;
        		o22cld_apparent_scene_pressure:units = "Pa" ;
        		o22cld_apparent_scene_pressure:long_name = "air_pressure_at_cloud_optical_centroid_assuming_completely_cloudy_sky" ;
        		o22cld_apparent_scene_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_apparent_scene_pressure:ancillary_variables = "o22cld_apparent_scene_pressure_precision" ;
        		o22cld_apparent_scene_pressure:_FillValue = 9.96921e+36f ;
        	float o22cld_apparent_scene_pressure_precision(time, scanline, ground_pixel) ;
        		o22cld_apparent_scene_pressure_precision:units = "Pa" ;
        		o22cld_apparent_scene_pressure_precision:long_name = "air_pressure_at_cloud_optical_centroid_assuming_completely_cloudy_sky standard_error" ;
        		o22cld_apparent_scene_pressure_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_apparent_scene_pressure_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_chi_square(time, scanline, ground_pixel) ;
        		o22cld_chi_square:units = "1" ;
        		o22cld_chi_square:long_name = "chi squared parameter of O2-O2 cloud fit" ;
        		o22cld_chi_square:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_chi_square:_FillValue = 9.96921e+36f ;
        	float o22cld_continuum_at_reference_wavelength(time, scanline, ground_pixel) ;
        		o22cld_continuum_at_reference_wavelength:units = "1" ;
        		o22cld_continuum_at_reference_wavelength:long_name = "continuum_reflectance_at_reference_wavelength" ;
        		o22cld_continuum_at_reference_wavelength:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_continuum_at_reference_wavelength:reference_wavelength = 475.f ;
        		o22cld_continuum_at_reference_wavelength:ancillary_variables = "o22cld_continuum_at_reference_wavelength_precision" ;
        		o22cld_continuum_at_reference_wavelength:_FillValue = 9.96921e+36f ;
        	float o22cld_continuum_at_reference_wavelength_precision(time, scanline, ground_pixel) ;
        		o22cld_continuum_at_reference_wavelength_precision:units = "1" ;
        		o22cld_continuum_at_reference_wavelength_precision:long_name = "continuum_reflectance_at_reference_wavelength standard_error" ;
        		o22cld_continuum_at_reference_wavelength_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_continuum_at_reference_wavelength_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_polynomial_coefficient(time, scanline, ground_pixel) ;
        		o22cld_polynomial_coefficient:units = "1" ;
        		o22cld_polynomial_coefficient:long_name = "first_order_background_polynomial_coefficient" ;
        		o22cld_polynomial_coefficient:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_polynomial_coefficient:reference_wavelength = 475.f ;
        		o22cld_polynomial_coefficient:ancillary_variables = "o22cld_polynomial_coefficient_precision" ;
        		o22cld_polynomial_coefficient:_FillValue = 9.96921e+36f ;
        	float o22cld_polynomial_coefficient_precision(time, scanline, ground_pixel) ;
        		o22cld_polynomial_coefficient_precision:units = "1" ;
        		o22cld_polynomial_coefficient_precision:long_name = "first_order_background_polynomial_coefficient standard_error" ;
        		o22cld_polynomial_coefficient_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_polynomial_coefficient_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_ring_coefficient(time, scanline, ground_pixel) ;
        		o22cld_ring_coefficient:units = "1" ;
        		o22cld_ring_coefficient:long_name = "ring_coefficient" ;
        		o22cld_ring_coefficient:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_ring_coefficient:ancillary_variables = "o22cld_ring_coefficient_precision" ;
        		o22cld_ring_coefficient:_FillValue = 9.96921e+36f ;
        	float o22cld_ring_coefficient_precision(time, scanline, ground_pixel) ;
        		o22cld_ring_coefficient_precision:units = "1" ;
        		o22cld_ring_coefficient_precision:long_name = "ring_coefficient standard_error" ;
        		o22cld_ring_coefficient_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_ring_coefficient_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_nitrogendioxide_slant_column_density(time, scanline, ground_pixel) ;
        		o22cld_nitrogendioxide_slant_column_density:units = "mol m-2" ;
        		o22cld_nitrogendioxide_slant_column_density:long_name = "slant_column_density_of_nitrogen_dioxide" ;
        		o22cld_nitrogendioxide_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_nitrogendioxide_slant_column_density:ancillary_variables = "o22cld_nitrogendioxide_slant_column_density_precision" ;
        		o22cld_nitrogendioxide_slant_column_density:_FillValue = 9.96921e+36f ;
        	float o22cld_nitrogendioxide_slant_column_density_precision(time, scanline, ground_pixel) ;
        		o22cld_nitrogendioxide_slant_column_density_precision:units = "mol m-2" ;
        		o22cld_nitrogendioxide_slant_column_density_precision:long_name = "slant_column_density_of_nitrogen_dioxide standard_error" ;
        		o22cld_nitrogendioxide_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_nitrogendioxide_slant_column_density_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_oxygen_oxygen_dimer_slant_column_density(time, scanline, ground_pixel) ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density:units = "mol2 m-5" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density:long_name = "slant_column_density_of_oxygen_cia" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density:ancillary_variables = "o22cld_oxygen_oxygen_dimer_slant_column_density_precision o22cld_oxygen_oxygen_dimer_slant_column_density_correction_factor" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density:_FillValue = 9.96921e+36f ;
        	float o22cld_oxygen_oxygen_dimer_slant_column_density_precision(time, scanline, ground_pixel) ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_precision:units = "mol2 m-5" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_precision:long_name = "slant_column_density_of_oxygen_cia standard_error" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_oxygen_oxygen_dimer_slant_column_density_correction_factor(time, scanline, ground_pixel) ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_correction_factor:units = "1" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_correction_factor:long_name = "O2-O2 slant column density temperature profile correction factor" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_correction_factor:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_oxygen_oxygen_dimer_slant_column_density_correction_factor:_FillValue = 9.96921e+36f ;
        	float o22cld_ozone_slant_column_density(time, scanline, ground_pixel) ;
        		o22cld_ozone_slant_column_density:units = "mol m-2" ;
        		o22cld_ozone_slant_column_density:long_name = "slant_column_density_of_ozone" ;
        		o22cld_ozone_slant_column_density:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_ozone_slant_column_density:ancillary_variables = "o22cld_ozone_slant_column_density_precision" ;
        		o22cld_ozone_slant_column_density:_FillValue = 9.96921e+36f ;
        	float o22cld_ozone_slant_column_density_precision(time, scanline, ground_pixel) ;
        		o22cld_ozone_slant_column_density_precision:units = "mol m-2" ;
        		o22cld_ozone_slant_column_density_precision:long_name = "slant_column_density_of_ozone standard_error" ;
        		o22cld_ozone_slant_column_density_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_ozone_slant_column_density_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_surface_albedo(time, scanline, ground_pixel) ;
        		o22cld_surface_albedo:units = "1" ;
        		o22cld_surface_albedo:standard_name = "surface_albedo" ;
        		o22cld_surface_albedo:long_name = "assumed surface albedo at 475 nm" ;
        		o22cld_surface_albedo:radiation_wavelength = 475.f ;
        		o22cld_surface_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_surface_albedo:_FillValue = 9.96921e+36f ;
        	float o22cld_wavelength_calibration_irradiance_offset(time, ground_pixel) ;
        		o22cld_wavelength_calibration_irradiance_offset:long_name = "wavelength offset" ;
        		o22cld_wavelength_calibration_irradiance_offset:units = "nm" ;
        		o22cld_wavelength_calibration_irradiance_offset:wavelength_fit_window_start = 460. ;
        		o22cld_wavelength_calibration_irradiance_offset:wavelength_fit_window_end = 490. ;
        		o22cld_wavelength_calibration_irradiance_offset:comment = "True wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
        		o22cld_wavelength_calibration_irradiance_offset:_FillValue = 9.96921e+36f ;
        	float o22cld_wavelength_calibration_irradiance_offset_precision(time, ground_pixel) ;
        		o22cld_wavelength_calibration_irradiance_offset_precision:long_name = "wavelength offset precision for the O2-O2 cloud parameters" ;
        		o22cld_wavelength_calibration_irradiance_offset_precision:units = "nm" ;
        		o22cld_wavelength_calibration_irradiance_offset_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_wavelength_calibration_irradiance_offset_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_wavelength_calibration_offset(time, scanline, ground_pixel) ;
        		o22cld_wavelength_calibration_offset:long_name = "wavelength offset" ;
        		o22cld_wavelength_calibration_offset:units = "nm" ;
        		o22cld_wavelength_calibration_offset:wavelength_fit_window_start = 460. ;
        		o22cld_wavelength_calibration_offset:wavelength_fit_window_end = 490. ;
        		o22cld_wavelength_calibration_offset:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_wavelength_calibration_offset:ancillary_variables = "o22cld_wavelength_calibration_offset_precision" ;
        		o22cld_wavelength_calibration_offset:comment = "True wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
        		o22cld_wavelength_calibration_offset:_FillValue = 9.96921e+36f ;
        	float o22cld_wavelength_calibration_offset_precision(time, scanline, ground_pixel) ;
        		o22cld_wavelength_calibration_offset_precision:long_name = "wavelength offset precision" ;
        		o22cld_wavelength_calibration_offset_precision:units = "nm" ;
        		o22cld_wavelength_calibration_offset_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_wavelength_calibration_offset_precision:_FillValue = 9.96921e+36f ;
        	float o22cld_wavelength_calibration_stretch(time, scanline, ground_pixel) ;
        		o22cld_wavelength_calibration_stretch:long_name = "wavelength stretch" ;
        		o22cld_wavelength_calibration_stretch:units = "1" ;
        		o22cld_wavelength_calibration_stretch:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_wavelength_calibration_stretch:ancillary_variables = "o22cld_wavelength_calibration_stretch_precision" ;
        		o22cld_wavelength_calibration_stretch:comment = "True wavelength = nominal wavelength + wavelength offset + wavelength stretch * scaled wavelength" ;
        		o22cld_wavelength_calibration_stretch:_FillValue = 9.96921e+36f ;
        	float o22cld_wavelength_calibration_stretch_precision(time, scanline, ground_pixel) ;
        		o22cld_wavelength_calibration_stretch_precision:long_name = "wavelength stretch precision" ;
        		o22cld_wavelength_calibration_stretch_precision:units = "1" ;
        		o22cld_wavelength_calibration_stretch_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		o22cld_wavelength_calibration_stretch_precision:_FillValue = 9.96921e+36f ;

        // group attributes:
        		:comment = "Cloud O2-O2 results" ;
        } // group O22CLD

      group: FRESCO {
        variables:
        	float fresco_cloud_fraction_crb(time, scanline, ground_pixel) ;
        		fresco_cloud_fraction_crb:units = "1" ;
        		fresco_cloud_fraction_crb:long_name = "effective_cloud_area_fraction_assuming_fixed_cloud_albedo" ;
        		fresco_cloud_fraction_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		fresco_cloud_fraction_crb:_FillValue = 9.96921e+36f ;
        	float fresco_cloud_pressure_crb(time, scanline, ground_pixel) ;
        		fresco_cloud_pressure_crb:units = "Pa" ;
        		fresco_cloud_pressure_crb:long_name = "air_pressure_at_cloud_optical_centroid" ;
        		fresco_cloud_pressure_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		fresco_cloud_pressure_crb:_FillValue = 9.96921e+36f ;
        	float fresco_scene_albedo(time, scanline, ground_pixel) ;
        		fresco_scene_albedo:units = "1" ;
        		fresco_scene_albedo:radiation_wavelength = 758.f ;
        		fresco_scene_albedo:long_name = "cloud_albedo_assuming_completely_cloudy_sky" ;
        		fresco_scene_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		fresco_scene_albedo:_FillValue = 9.96921e+36f ;
        	float fresco_apparent_scene_pressure(time, scanline, ground_pixel) ;
        		fresco_apparent_scene_pressure:units = "Pa" ;
        		fresco_apparent_scene_pressure:long_name = "air_pressure_at_cloud_optical_centroid_assuming_completely_cloudy_sky" ;
        		fresco_apparent_scene_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
        		fresco_apparent_scene_pressure:_FillValue = 9.96921e+36f ;
        	float fresco_cloud_albedo_crb(time, scanline, ground_pixel) ;
        		fresco_cloud_albedo_crb:units = "1" ;
        		fresco_cloud_albedo_crb:standard_name = "cloud_albedo" ;
        		fresco_cloud_albedo_crb:long_name = "cloud albedo" ;
        		fresco_cloud_albedo_crb:coordinates = "longitude latitude" ;
        		fresco_cloud_albedo_crb:ancillary_variables = "cloud_albedo_precision" ;
        		fresco_cloud_albedo_crb:_FillValue = 9.96921e+36f ;
        	float fresco_surface_albedo(time, scanline, ground_pixel) ;
        		fresco_surface_albedo:units = "1" ;
        		fresco_surface_albedo:standard_name = "surface_albedo" ;
        		fresco_surface_albedo:long_name = "assumed surface albedo at 758 nm" ;
        		fresco_surface_albedo:radiation_wavelength = 758.f ;
        		fresco_surface_albedo:coordinates = "longitude latitude" ;
        		fresco_surface_albedo:_FillValue = 9.96921e+36f ;

        // group attributes:
        		:comment = "Remapped FRESCO results" ;
        } // group FRESCO
      } // group DETAILED_RESULTS

    group: INPUT_DATA {
      variables:
      	float surface_altitude(time, scanline, ground_pixel) ;
      		surface_altitude:long_name = "Surface altitude" ;
      		surface_altitude:standard_name = "surface_altitude" ;
      		surface_altitude:units = "m" ;
      		surface_altitude:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude:comment = "The mean of the sub-pixels of the surface altitudewithin the approximate field of view, based on the GMTED2010 surface elevation database" ;
      		surface_altitude:_FillValue = 9.96921e+36f ;
      	float surface_altitude_precision(time, scanline, ground_pixel) ;
      		surface_altitude_precision:long_name = "surface altitude precision" ;
      		surface_altitude_precision:standard_name = "surface_altitude standard_error" ;
      		surface_altitude_precision:units = "m" ;
      		surface_altitude_precision:standard_error_multiplier = 1.f ;
      		surface_altitude_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude_precision:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude_precision:comment = "The standard deviation of sub-pixels used in calculating the mean surface altitude, based on the GMTED2010 surface elevation database" ;
      		surface_altitude_precision:_FillValue = 9.96921e+36f ;
      	ubyte surface_classification(time, scanline, ground_pixel) ;
      		surface_classification:long_name = "Land-water mask and surface classification based on a static database" ;
      		surface_classification:comment = "Flag indicating land/water and further surface classifications for the ground pixel" ;
      		surface_classification:source = "USGS (https://lta.cr.usgs.gov/GLCC) and NASA SDP toolkit (http://newsroom.gsfc.nasa.gov/sdptoolkit/toolkit.html)" ;
      		surface_classification:flag_meanings = "land water some_water coast value_covers_majority_of_pixel water+shallow_ocean water+shallow_inland_water water+ocean_coastline-lake_shoreline water+intermittent_water water+deep_inland_water water+continental_shelf_ocean water+deep_ocean land+urban_and_built-up_land land+dryland_cropland_and_pasture land+irrigated_cropland_and_pasture land+mixed_dryland-irrigated_cropland_and_pasture land+cropland-grassland_mosaic land+cropland-woodland_mosaic land+grassland land+shrubland land+mixed_shrubland-grassland land+savanna land+deciduous_broadleaf_forest land+deciduous_needleleaf_forest land+evergreen_broadleaf_forest land+evergreen_needleleaf_forest land+mixed_forest land+herbaceous_wetland land+wooded_wetland land+barren_or_sparsely_vegetated land+herbaceous_tundra land+wooded_tundra land+mixed_tundra land+bare_ground_tundra land+snow_or_ice" ;
      		surface_classification:flag_values = 0UB, 1UB, 2UB, 3UB, 4UB, 9UB, 17UB, 25UB, 33UB, 41UB, 49UB, 57UB, 8UB, 16UB, 24UB, 32UB, 40UB, 48UB, 56UB, 64UB, 72UB, 80UB, 88UB, 96UB, 104UB, 112UB, 120UB, 128UB, 136UB, 144UB, 152UB, 160UB, 168UB, 176UB, 184UB ;
      		surface_classification:flag_masks = 3UB, 3UB, 3UB, 3UB, 4UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB ;
      		surface_classification:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_classification:_FillValue = 255UB ;
      	int instrument_configuration_identifier(time, scanline) ;
      		instrument_configuration_identifier:long_name = "IcID" ;
      		instrument_configuration_identifier:comment = "The Instrument Configuration ID defines the type of measurement and its purpose. The number of instrument configuration IDs will increase over the mission as new types of measurements are created and used" ;
      		instrument_configuration_identifier:_FillValue = -2147483647 ;
      	short instrument_configuration_version(time, scanline) ;
      		instrument_configuration_version:long_name = "IcVersion" ;
      		instrument_configuration_version:comment = "Version of the instrument_configuration_identifier" ;
      		instrument_configuration_version:_FillValue = -32767s ;
      	float scaled_small_pixel_variance(time, scanline, ground_pixel) ;
      		scaled_small_pixel_variance:long_name = "scaled small pixel variance" ;
      		scaled_small_pixel_variance:units = "1" ;
      		scaled_small_pixel_variance:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		scaled_small_pixel_variance:comment = "The scaled variance of the reflectances of the small pixels" ;
      		scaled_small_pixel_variance:radiation_wavelength = 460.f ;
      		scaled_small_pixel_variance:_FillValue = 9.96921e+36f ;
      	float eastward_wind(time, scanline, ground_pixel) ;
      		eastward_wind:standard_name = "eastward_wind" ;
      		eastward_wind:long_name = "Eastward wind from ECMWF at 10 meter height level" ;
      		eastward_wind:units = "m s-1" ;
      		eastward_wind:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		eastward_wind:ancillary_variables = "northward_wind" ;
      		eastward_wind:_FillValue = 9.96921e+36f ;
      	float northward_wind(time, scanline, ground_pixel) ;
      		northward_wind:standard_name = "northward_wind" ;
      		northward_wind:long_name = "Northward wind from ECMWF at 10 meter height level" ;
      		northward_wind:units = "m s-1" ;
      		northward_wind:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		northward_wind:ancillary_variables = "eastward_wind" ;
      		northward_wind:_FillValue = 9.96921e+36f ;
      	float surface_pressure(time, scanline, ground_pixel) ;
      		surface_pressure:units = "Pa" ;
      		surface_pressure:standard_name = "surface_air_pressure" ;
      		surface_pressure:long_name = "Surface pressure" ;
      		surface_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_pressure:_FillValue = 9.96921e+36f ;
      	float surface_albedo_nitrogendioxide_window(time, scanline, ground_pixel) ;
      		surface_albedo_nitrogendioxide_window:units = "1" ;
      		surface_albedo_nitrogendioxide_window:standard_name = "surface_albedo" ;
      		surface_albedo_nitrogendioxide_window:long_name = "Surface albedo in the NO2 fit window" ;
      		surface_albedo_nitrogendioxide_window:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_albedo_nitrogendioxide_window:_FillValue = 9.96921e+36f ;
      	float surface_albedo(time, scanline, ground_pixel) ;
      		surface_albedo:units = "1" ;
      		surface_albedo:standard_name = "surface_albedo" ;
      		surface_albedo:long_name = "Surface albedo in the cloud product" ;
      		surface_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_albedo:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/cloud_selection_flag" ;
      		surface_albedo:_FillValue = 9.96921e+36f ;
      	float cloud_pressure_crb(time, scanline, ground_pixel) ;
      		cloud_pressure_crb:units = "Pa" ;
      		cloud_pressure_crb:proposed_standard_name = "air_pressure_at_cloud_optical_centroid" ;
      		cloud_pressure_crb:long_name = "Cloud optical centroid pressure" ;
      		cloud_pressure_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_pressure_crb:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/cloud_selection_flag" ;
      		cloud_pressure_crb:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_crb(time, scanline, ground_pixel) ;
      		cloud_fraction_crb:units = "1" ;
      		cloud_fraction_crb:proposed_standard_name = "effective_cloud_area_fraction_assuming_fixed_cloud_albedo" ;
      		cloud_fraction_crb:long_name = "Effective cloud fraction from the cloud product" ;
      		cloud_fraction_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_crb:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/cloud_selection_flag" ;
      		cloud_fraction_crb:_FillValue = 9.96921e+36f ;
      	float cloud_albedo_crb(time, scanline, ground_pixel) ;
      		cloud_albedo_crb:units = "1" ;
      		cloud_albedo_crb:standard_name = "cloud_albedo" ;
      		cloud_albedo_crb:long_name = "Cloud albedo in the cloud product" ;
      		cloud_albedo_crb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_albedo_crb:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/cloud_selection_flag" ;
      		cloud_albedo_crb:_FillValue = 9.96921e+36f ;
      	float scene_albedo(time, scanline, ground_pixel) ;
      		scene_albedo:units = "1" ;
      		scene_albedo:proposed_standard_name = "cloud_albedo_assuming_completely_cloudy_sky" ;
      		scene_albedo:long_name = "Scene albedo in the cloud product" ;
      		scene_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		scene_albedo:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/cloud_selection_flag" ;
      		scene_albedo:_FillValue = 9.96921e+36f ;
      	float apparent_scene_pressure(time, scanline, ground_pixel) ;
      		apparent_scene_pressure:units = "Pa" ;
      		apparent_scene_pressure:proposed_standard_name = "air_pressure_at_cloud_optical_centroid_assuming_completely_cloudy_sky" ;
      		apparent_scene_pressure:long_name = "Scene pressure from the cloud product" ;
      		apparent_scene_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		apparent_scene_pressure:ancillary_variables = "/PRODUCT/SUPPORT_DATA/DETAILED_RESULTS/cloud_selection_flag" ;
      		apparent_scene_pressure:_FillValue = 9.96921e+36f ;
      	ubyte snow_ice_flag(time, scanline, ground_pixel) ;
      		snow_ice_flag:long_name = "Snow-ice mask" ;
      		snow_ice_flag:_FillValue = 254UB ;
      		snow_ice_flag:comment = "Flag indicating snow/ice at center of ground pixel" ;
      		snow_ice_flag:source = "ECMWF" ;
      		snow_ice_flag:flag_meanings = "snow-free_land sea_ice_1_percent sea_ice_2_percent sea_ice_3_percent sea_ice_4_percent sea_ice_5_percent sea_ice_6_percent sea_ice_7_percent sea_ice_8_percent sea_ice_9_percent sea_ice_10_percent sea_ice_11_percent sea_ice_12_percent sea_ice_13_percent sea_ice_14_percent sea_ice_15_percent sea_ice_16_percent sea_ice_17_percent sea_ice_18_percent sea_ice_19_percent sea_ice_20_percent sea_ice_21_percent sea_ice_22_percent sea_ice_23_percent sea_ice_24_percent sea_ice_25_percent sea_ice_26_percent sea_ice_27_percent sea_ice_28_percent sea_ice_29_percent sea_ice_30_percent sea_ice_31_percent sea_ice_32_percent sea_ice_33_percent sea_ice_34_percent sea_ice_35_percent sea_ice_36_percent sea_ice_37_percent sea_ice_38_percent sea_ice_39_percent sea_ice_40_percent sea_ice_41_percent sea_ice_42_percent sea_ice_43_percent sea_ice_44_percent sea_ice_45_percent sea_ice_46_percent sea_ice_47_percent sea_ice_48_percent sea_ice_49_percent sea_ice_50_percent sea_ice_51_percent sea_ice_52_percent sea_ice_53_percent sea_ice_54_percent sea_ice_55_percent sea_ice_56_percent sea_ice_57_percent sea_ice_58_percent sea_ice_59_percent sea_ice_60_percent sea_ice_61_percent sea_ice_62_percent sea_ice_63_percent sea_ice_64_percent sea_ice_65_percent sea_ice_66_percent sea_ice_67_percent sea_ice_68_percent sea_ice_69_percent sea_ice_70_percent sea_ice_71_percent sea_ice_72_percent sea_ice_73_percent sea_ice_74_percent sea_ice_75_percent sea_ice_76_percent sea_ice_77_percent sea_ice_78_percent sea_ice_79_percent sea_ice_80_percent sea_ice_81_percent sea_ice_82_percent sea_ice_83_percent sea_ice_84_percent sea_ice_85_percent sea_ice_86_percent sea_ice_87_percent sea_ice_88_percent sea_ice_89_percent sea_ice_90_percent sea_ice_91_percent sea_ice_92_percent sea_ice_93_percent sea_ice_94_percent sea_ice_95_percent sea_ice_96_percent sea_ice_97_percent sea_ice_98_percent sea_ice_99_percent sea_ice_100_percent permanent_ice snow mixed_pixels_at_coastlines suspect_ice_value corners ocean" ;
      		snow_ice_flag:flag_values = 0UB, 1UB, 2UB, 3UB, 4UB, 5UB, 6UB, 7UB, 8UB, 9UB, 10UB, 11UB, 12UB, 13UB, 14UB, 15UB, 16UB, 17UB, 18UB, 19UB, 20UB, 21UB, 22UB, 23UB, 24UB, 25UB, 26UB, 27UB, 28UB, 29UB, 30UB, 31UB, 32UB, 33UB, 34UB, 35UB, 36UB, 37UB, 38UB, 39UB, 40UB, 41UB, 42UB, 43UB, 44UB, 45UB, 46UB, 47UB, 48UB, 49UB, 50UB, 51UB, 52UB, 53UB, 54UB, 55UB, 56UB, 57UB, 58UB, 59UB, 60UB, 61UB, 62UB, 63UB, 64UB, 65UB, 66UB, 67UB, 68UB, 69UB, 70UB, 71UB, 72UB, 73UB, 74UB, 75UB, 76UB, 77UB, 78UB, 79UB, 80UB, 81UB, 82UB, 83UB, 84UB, 85UB, 86UB, 87UB, 88UB, 89UB, 90UB, 91UB, 92UB, 93UB, 94UB, 95UB, 96UB, 97UB, 98UB, 99UB, 100UB, 101UB, 103UB, 252UB, 253UB, 254UB, 255UB ;
      		snow_ice_flag:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float aerosol_index_354_388(time, scanline, ground_pixel) ;
      		aerosol_index_354_388:units = "1" ;
      		aerosol_index_354_388:long_name = "Absorbing aerosol index from the TROPOMI AAI product" ;
      		aerosol_index_354_388:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_index_354_388:_FillValue = 9.96921e+36f ;
      } // group INPUT_DATA
    } // group SUPPORT_DATA
  } // group PRODUCT

group: METADATA {

  group: QA_STATISTICS {
    dimensions:
    	vertices = 2 ;
    	nitrogendioxide_tropospheric_column_histogram_axis = 100 ;
    	nitrogendioxide_tropospheric_column_pdf_axis = 400 ;
    	nitrogendioxide_stratospheric_column_histogram_axis = 100 ;
    	nitrogendioxide_stratospheric_column_pdf_axis = 400 ;
    	nitrogendioxide_total_column_histogram_axis = 100 ;
    	nitrogendioxide_total_column_pdf_axis = 400 ;
    variables:
    	float nitrogendioxide_stratospheric_column_histogram_axis(nitrogendioxide_stratospheric_column_histogram_axis) ;
    		nitrogendioxide_stratospheric_column_histogram_axis:units = "mol m-2" ;
    		nitrogendioxide_stratospheric_column_histogram_axis:comment = "Histogram of the stratospheric NO2 vertical column" ;
    		nitrogendioxide_stratospheric_column_histogram_axis:long_name = "Histogram of the stratospheric NO2 vertical column" ;
    		nitrogendioxide_stratospheric_column_histogram_axis:bounds = "nitrogendioxide_stratospheric_column_histogram_bounds" ;
    		nitrogendioxide_stratospheric_column_histogram_axis:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_stratospheric_column_pdf_axis(nitrogendioxide_stratospheric_column_pdf_axis) ;
    		nitrogendioxide_stratospheric_column_pdf_axis:units = "mol m-2" ;
    		nitrogendioxide_stratospheric_column_pdf_axis:comment = "Probability density function of the stratospheric NO2 vertical column" ;
    		nitrogendioxide_stratospheric_column_pdf_axis:long_name = "Probability density function of the stratospheric NO2 vertical column" ;
    		nitrogendioxide_stratospheric_column_pdf_axis:bounds = "aerosol_nitrogendioxide_stratospheric_column_pdf_bounds" ;
    		nitrogendioxide_stratospheric_column_pdf_axis:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_stratospheric_column_histogram_bounds(nitrogendioxide_stratospheric_column_histogram_axis, vertices) ;
    		nitrogendioxide_stratospheric_column_histogram_bounds:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_stratospheric_column_pdf_bounds(nitrogendioxide_stratospheric_column_pdf_axis, vertices) ;
    		nitrogendioxide_stratospheric_column_pdf_bounds:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_tropospheric_column_histogram_axis(nitrogendioxide_tropospheric_column_histogram_axis) ;
    		nitrogendioxide_tropospheric_column_histogram_axis:units = "mol m-2" ;
    		nitrogendioxide_tropospheric_column_histogram_axis:comment = "Histogram of the tropospheric NO2 vertical column" ;
    		nitrogendioxide_tropospheric_column_histogram_axis:long_name = "Histogram of the tropospheric NO2 vertical column" ;
    		nitrogendioxide_tropospheric_column_histogram_axis:bounds = "nitrogendioxide_tropospheric_column_histogram_bounds" ;
    		nitrogendioxide_tropospheric_column_histogram_axis:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_tropospheric_column_pdf_axis(nitrogendioxide_tropospheric_column_pdf_axis) ;
    		nitrogendioxide_tropospheric_column_pdf_axis:units = "mol m-2" ;
    		nitrogendioxide_tropospheric_column_pdf_axis:comment = "Probability density function of the tropospheric NO2 vertical column" ;
    		nitrogendioxide_tropospheric_column_pdf_axis:long_name = "Probability density function of the tropospheric NO2 vertical column" ;
    		nitrogendioxide_tropospheric_column_pdf_axis:bounds = "nitrogendioxide_tropospheric_column_pdf_bounds" ;
    		nitrogendioxide_tropospheric_column_pdf_axis:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_tropospheric_column_histogram_bounds(nitrogendioxide_tropospheric_column_histogram_axis, vertices) ;
    		nitrogendioxide_tropospheric_column_histogram_bounds:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_tropospheric_column_pdf_bounds(nitrogendioxide_tropospheric_column_pdf_axis, vertices) ;
    		nitrogendioxide_tropospheric_column_pdf_bounds:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_total_column_histogram_axis(nitrogendioxide_total_column_histogram_axis) ;
    		nitrogendioxide_total_column_histogram_axis:units = "mol m-2" ;
    		nitrogendioxide_total_column_histogram_axis:comment = "Histogram of the total NO2 vertical column" ;
    		nitrogendioxide_total_column_histogram_axis:long_name = "Histogram of the total NO2 vertical column" ;
    		nitrogendioxide_total_column_histogram_axis:bounds = "nitrogendioxide_total_column_histogram_bounds" ;
    		nitrogendioxide_total_column_histogram_axis:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_total_column_pdf_axis(nitrogendioxide_total_column_pdf_axis) ;
    		nitrogendioxide_total_column_pdf_axis:units = "mol m-2" ;
    		nitrogendioxide_total_column_pdf_axis:comment = "Probability density function of the total NO2 vertical column" ;
    		nitrogendioxide_total_column_pdf_axis:long_name = "Probability density function of the total NO2 vertical column" ;
    		nitrogendioxide_total_column_pdf_axis:bounds = "nitrogendioxide_total_column_pdf_bounds" ;
    		nitrogendioxide_total_column_pdf_axis:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_total_column_histogram_bounds(nitrogendioxide_total_column_histogram_axis, vertices) ;
    		nitrogendioxide_total_column_histogram_bounds:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_total_column_pdf_bounds(nitrogendioxide_total_column_pdf_axis, vertices) ;
    		nitrogendioxide_total_column_pdf_bounds:_FillValue = 9.96921e+36f ;
    	int nitrogendioxide_tropospheric_column_histogram(nitrogendioxide_tropospheric_column_histogram_axis) ;
    		nitrogendioxide_tropospheric_column_histogram:comment = "Histogram of the tropospheric NO2 vertical column in the current granule" ;
    		nitrogendioxide_tropospheric_column_histogram:number_of_overflow_values = 46 ;
    		nitrogendioxide_tropospheric_column_histogram:number_of_underflow_values = 90461 ;
    		nitrogendioxide_tropospheric_column_histogram:_FillValue = -2147483647 ;
    	int nitrogendioxide_stratospheric_column_histogram(nitrogendioxide_stratospheric_column_histogram_axis) ;
    		nitrogendioxide_stratospheric_column_histogram:comment = "Histogram of the stratospheric NO2 vertical column in the current granule" ;
    		nitrogendioxide_stratospheric_column_histogram:number_of_overflow_values = 0 ;
    		nitrogendioxide_stratospheric_column_histogram:number_of_underflow_values = 0 ;
    		nitrogendioxide_stratospheric_column_histogram:_FillValue = -2147483647 ;
    	int nitrogendioxide_total_column_histogram(nitrogendioxide_total_column_histogram_axis) ;
    		nitrogendioxide_total_column_histogram:comment = "Histogram of the total NO2 vertical column in the current granule" ;
    		nitrogendioxide_total_column_histogram:number_of_overflow_values = 0 ;
    		nitrogendioxide_total_column_histogram:number_of_underflow_values = 0 ;
    		nitrogendioxide_total_column_histogram:_FillValue = -2147483647 ;
    	float nitrogendioxide_tropospheric_column_pdf(nitrogendioxide_tropospheric_column_pdf_axis) ;
    		nitrogendioxide_tropospheric_column_pdf:comment = "Probability density function of the tropospheric NO2 vertical column in the current granule" ;
    		nitrogendioxide_tropospheric_column_pdf:geolocation_sampling_total = 52630.21f ;
    		nitrogendioxide_tropospheric_column_pdf:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_stratospheric_column_pdf(nitrogendioxide_stratospheric_column_pdf_axis) ;
    		nitrogendioxide_stratospheric_column_pdf:comment = "Probability density function of the stratospheric NO2 vertical column in the current granule" ;
    		nitrogendioxide_stratospheric_column_pdf:geolocation_sampling_total = 113866.7f ;
    		nitrogendioxide_stratospheric_column_pdf:_FillValue = 9.96921e+36f ;
    	float nitrogendioxide_total_column_pdf(nitrogendioxide_total_column_pdf_axis) ;
    		nitrogendioxide_total_column_pdf:comment = "Probability density function of the total NO2 vertical column in the current granule" ;
    		nitrogendioxide_total_column_pdf:geolocation_sampling_total = 113866.7f ;
    		nitrogendioxide_total_column_pdf:_FillValue = 9.96921e+36f ;

    // group attributes:
    		:number_of_groundpixels = 167400 ;
    		:number_of_processed_pixels = 167400 ;
    		:number_of_successfully_processed_pixels = 163287 ;
    		:number_of_rejected_pixels_not_enough_spectrum = 0 ;
    		:number_of_failed_retrievals = 4113 ;
    		:number_of_ground_pixels_with_warnings = 131843 ;
    		:number_of_missing_scanlines = 0 ;
    		:number_of_radiance_missing_occurrences = 0 ;
    		:number_of_irradiance_missing_occurrences = 0 ;
    		:number_of_input_spectrum_missing_occurrences = 0 ;
    		:number_of_reflectance_range_error_occurrences = 0 ;
    		:number_of_ler_range_error_occurrences = 0 ;
    		:number_of_snr_range_error_occurrences = 0 ;
    		:number_of_sza_range_error_occurrences = 0 ;
    		:number_of_vza_range_error_occurrences = 0 ;
    		:number_of_lut_range_error_occurrences = 0 ;
    		:number_of_ozone_range_error_occurrences = 0 ;
    		:number_of_wavelength_offset_error_occurrences = 0 ;
    		:number_of_initialization_error_occurrences = 0 ;
    		:number_of_memory_error_occurrences = 0 ;
    		:number_of_assertion_error_occurrences = 0 ;
    		:number_of_io_error_occurrences = 0 ;
    		:number_of_numerical_error_occurrences = 0 ;
    		:number_of_lut_error_occurrences = 0 ;
    		:number_of_ISRF_error_occurrences = 0 ;
    		:number_of_convergence_error_occurrences = 0 ;
    		:number_of_cloud_filter_convergence_error_occurrences = 0 ;
    		:number_of_max_iteration_convergence_error_occurrences = 0 ;
    		:number_of_aot_lower_boundary_convergence_error_occurrences = 0 ;
    		:number_of_other_boundary_convergence_error_occurrences = 0 ;
    		:number_of_geolocation_error_occurrences = 0 ;
    		:number_of_ch4_noscat_zero_error_occurrences = 0 ;
    		:number_of_h2o_noscat_zero_error_occurrences = 0 ;
    		:number_of_max_optical_thickness_error_occurrences = 0 ;
    		:number_of_aerosol_boundary_error_occurrences = 0 ;
    		:number_of_boundary_hit_error_occurrences = 0 ;
    		:number_of_chi2_error_occurrences = 0 ;
    		:number_of_svd_error_occurrences = 0 ;
    		:number_of_dfs_error_occurrences = 0 ;
    		:number_of_radiative_transfer_error_occurrences = 0 ;
    		:number_of_optimal_estimation_error_occurrences = 0 ;
    		:number_of_profile_error_occurrences = 0 ;
    		:number_of_cloud_error_occurrences = 4099 ;
    		:number_of_model_error_occurrences = 0 ;
    		:number_of_number_of_input_data_points_too_low_error_occurrences = 0 ;
    		:number_of_cloud_pressure_spread_too_low_error_occurrences = 0 ;
    		:number_of_cloud_too_low_level_error_occurrences = 0 ;
    		:number_of_generic_range_error_occurrences = 14 ;
    		:number_of_generic_exception_occurrences = 0 ;
    		:number_of_input_spectrum_alignment_error_occurrences = 0 ;
    		:number_of_abort_error_occurrences = 0 ;
    		:number_of_wrong_input_type_error_occurrences = 0 ;
    		:number_of_wavelength_calibration_error_occurrences = 0 ;
    		:number_of_coregistration_error_occurrences = 0 ;
    		:number_of_slant_column_density_error_occurrences = 0 ;
    		:number_of_airmass_factor_error_occurrences = 0 ;
    		:number_of_vertical_column_density_error_occurrences = 0 ;
    		:number_of_signal_to_noise_ratio_error_occurrences = 0 ;
    		:number_of_configuration_error_occurrences = 0 ;
    		:number_of_key_error_occurrences = 0 ;
    		:number_of_saturation_error_occurrences = 0 ;
    		:number_of_max_num_outlier_exceeded_error_occurrences = 0 ;
    		:number_of_solar_eclipse_filter_occurrences = 0 ;
    		:number_of_cloud_filter_occurrences = 0 ;
    		:number_of_altitude_consistency_filter_occurrences = 0 ;
    		:number_of_altitude_roughness_filter_occurrences = 0 ;
    		:number_of_sun_glint_filter_occurrences = 0 ;
    		:number_of_mixed_surface_type_filter_occurrences = 0 ;
    		:number_of_snow_ice_filter_occurrences = 0 ;
    		:number_of_aai_filter_occurrences = 0 ;
    		:number_of_cloud_fraction_fresco_filter_occurrences = 0 ;
    		:number_of_aai_scene_albedo_filter_occurrences = 0 ;
    		:number_of_small_pixel_radiance_std_filter_occurrences = 0 ;
    		:number_of_cloud_fraction_viirs_filter_occurrences = 0 ;
    		:number_of_cirrus_reflectance_viirs_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ifov_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofova_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofovb_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofovc_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ifov_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofova_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofovb_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofovc_filter_occurrences = 0 ;
    		:number_of_refl_cirrus_viirs_swir_filter_occurrences = 0 ;
    		:number_of_refl_cirrus_viirs_nir_filter_occurrences = 0 ;
    		:number_of_diff_refl_cirrus_viirs_filter_occurrences = 0 ;
    		:number_of_ch4_noscat_ratio_filter_occurrences = 0 ;
    		:number_of_ch4_noscat_ratio_std_filter_occurrences = 0 ;
    		:number_of_h2o_noscat_ratio_filter_occurrences = 0 ;
    		:number_of_h2o_noscat_ratio_std_filter_occurrences = 0 ;
    		:number_of_diff_psurf_fresco_ecmwf_filter_occurrences = 0 ;
    		:number_of_psurf_fresco_stdv_filter_occurrences = 0 ;
    		:number_of_ocean_filter_occurrences = 0 ;
    		:number_of_time_range_filter_occurrences = 0 ;
    		:number_of_pixel_or_scanline_index_filter_occurrences = 0 ;
    		:number_of_geographic_region_filter_occurrences = 0 ;
    		:number_of_internal_cloud_mask_filter_occurrences = 0 ;
    		:number_of_input_spectrum_warning_occurrences = 0 ;
    		:number_of_wavelength_calibration_warning_occurrences = 0 ;
    		:number_of_extrapolation_warning_occurrences = 0 ;
    		:number_of_sun_glint_warning_occurrences = 0 ;
    		:number_of_south_atlantic_anomaly_warning_occurrences = 0 ;
    		:number_of_sun_glint_correction_occurrences = 0 ;
    		:number_of_snow_ice_warning_occurrences = 119267 ;
    		:number_of_cloud_warning_occurrences = 0 ;
    		:number_of_AAI_warning_occurrences = 0 ;
    		:number_of_pixel_level_input_data_missing_occurrences = 18074 ;
    		:number_of_data_range_warning_occurrences = 0 ;
    		:number_of_low_cloud_fraction_warning_occurrences = 0 ;
    		:number_of_altitude_consistency_warning_occurrences = 0 ;
    		:number_of_signal_to_noise_ratio_warning_occurrences = 0 ;
    		:number_of_deconvolution_warning_occurrences = 0 ;
    		:number_of_so2_volcanic_origin_likely_warning_occurrences = 0 ;
    		:number_of_so2_volcanic_origin_certain_warning_occurrences = 0 ;
    		:number_of_interpolation_warning_occurrences = 0 ;
    		:number_of_saturation_warning_occurrences = 0 ;
    		:number_of_high_sza_warning_occurrences = 0 ;
    		:number_of_cloud_retrieval_warning_occurrences = 0 ;
    		:number_of_cloud_inhomogeneity_warning_occurrences = 0 ;
    		:number_of_thermal_instability_warning_occurrences = 0 ;
    		:global_processing_warnings = "None" ;
    		:time_for_algorithm_initialization = 97.764832 ;
    		:time_for_processing = 36.581845 ;
    		:time_per_pixel = 0.00557704501276885 ;
    		:time_standard_deviation_per_pixel = 1.00967782789192e-05 ;
    } // group QA_STATISTICS

  group: ALGORITHM_SETTINGS {

    // group attributes:
    		:CLDDOAS.NO2.output.name = "nitrogendioxide" ;
    		:CLDDOAS.O2O2.output.name = "oxygen_oxygen_dimer" ;
    		:CLDDOAS.O3.output.name = "ozone" ;
    		:CLDDOAS.background_offset.polynomial_order = "1" ;
    		:CLDDOAS.convergence_threshold = "1.0" ;
    		:CLDDOAS.filter_outliers = "true" ;
    		:CLDDOAS.filter_outliers_fraction = "0.0" ;
    		:CLDDOAS.filter_outliers_maximum_number_allowed_outliers = "5" ;
    		:CLDDOAS.filter_outliers_threshold = "3.0" ;
    		:CLDDOAS.include_offset = "false" ;
    		:CLDDOAS.include_ring = "true" ;
    		:CLDDOAS.initial_guess.NO2 = "1.8e-4" ;
    		:CLDDOAS.initial_guess.O2O2 = "8.0e+5" ;
    		:CLDDOAS.initial_guess.O3 = "3.6e-1" ;
    		:CLDDOAS.initial_guess.a0 = "1.0" ;
    		:CLDDOAS.initial_guess.a1 = "0.125" ;
    		:CLDDOAS.initial_guess.ring = "0.06" ;
    		:CLDDOAS.intensity_offset_scalefactor = "1.0" ;
    		:CLDDOAS.max_iterations = "15" ;
    		:CLDDOAS.output.prefix = "o22cld_" ;
    		:CLDDOAS.polynomial_order = "1" ;
    		:CLDDOAS.scale_precision_with_chisq = "true" ;
    		:CLDDOAS.sigma.NO2 = "1.0e-2" ;
    		:CLDDOAS.sigma.O2O2 = "2.0e+6" ;
    		:CLDDOAS.sigma.O3 = "5.0e0" ;
    		:CLDDOAS.sigma.a0 = "1.0" ;
    		:CLDDOAS.sigma.a1 = "0.125" ;
    		:CLDDOAS.sigma.ring = "0.2" ;
    		:CLDDOAS.species = "O2O2, NO2, O3" ;
    		:CLDDOAS.wavelength_end = "490.0" ;
    		:CLDDOAS.wavelength_start = "460.0" ;
    		:CLDDOAS.write_diagnostic_output = "false" ;
    		:NO2DOAS.H2O_liquid.output.name = "water_liquid" ;
    		:NO2DOAS.H2O_vapor.output.name = "water" ;
    		:NO2DOAS.NO2.output.name = "nitrogendioxide" ;
    		:NO2DOAS.NO2.reference_temperature = "-1.0" ;
    		:NO2DOAS.O2O2.output.name = "oxygen_oxygen_dimer" ;
    		:NO2DOAS.O3.output.name = "ozone" ;
    		:NO2DOAS.O3.reference_temperature = "-1.0" ;
    		:NO2DOAS.background_offset.polynomial_order = "1" ;
    		:NO2DOAS.convergence_threshold = "0.99" ;
    		:NO2DOAS.filter_outliers = "true" ;
    		:NO2DOAS.filter_outliers_fraction = "0.0" ;
    		:NO2DOAS.filter_outliers_maximum_number_allowed_outliers = "10" ;
    		:NO2DOAS.filter_outliers_threshold = "3.0" ;
    		:NO2DOAS.include_offset = "false" ;
    		:NO2DOAS.include_ring = "true" ;
    		:NO2DOAS.initial_guess.H2O_liquid = "0.0" ;
    		:NO2DOAS.initial_guess.H2O_vapor = "1.5e+3" ;
    		:NO2DOAS.initial_guess.NO2 = "1.2e-5" ;
    		:NO2DOAS.initial_guess.O2O2 = "8.0e+5" ;
    		:NO2DOAS.initial_guess.O3 = "3.6e-1" ;
    		:NO2DOAS.initial_guess.a0 = "1.0" ;
    		:NO2DOAS.initial_guess.a1 = "0.125" ;
    		:NO2DOAS.initial_guess.a2 = "0.015625" ;
    		:NO2DOAS.initial_guess.a3 = "0.015625" ;
    		:NO2DOAS.initial_guess.a4 = "0.015625" ;
    		:NO2DOAS.initial_guess.a5 = "0.015625" ;
    		:NO2DOAS.initial_guess.c0 = "1.0" ;
    		:NO2DOAS.initial_guess.c1 = "0.125" ;
    		:NO2DOAS.initial_guess.c2 = "0.015625" ;
    		:NO2DOAS.initial_guess.c3 = "0.015625" ;
    		:NO2DOAS.initial_guess.ring = "0.06" ;
    		:NO2DOAS.intensity_offset_scalefactor = "1.0" ;
    		:NO2DOAS.max_iterations = "20" ;
    		:NO2DOAS.polynomial_order = "5" ;
    		:NO2DOAS.reference_cross_sections_key = "REF_XS_NO2" ;
    		:NO2DOAS.scale_precision_with_chisq = "true" ;
    		:NO2DOAS.sigma.H2O_liquid = "20.0" ;
    		:NO2DOAS.sigma.H2O_vapor = "1.0e+4" ;
    		:NO2DOAS.sigma.NO2 = "1.0e-2" ;
    		:NO2DOAS.sigma.O2O2 = "2.0e+6" ;
    		:NO2DOAS.sigma.O3 = "5.0e0" ;
    		:NO2DOAS.sigma.a0 = "1.0" ;
    		:NO2DOAS.sigma.a1 = "0.125" ;
    		:NO2DOAS.sigma.a2 = "0.015625" ;
    		:NO2DOAS.sigma.a3 = "0.015625" ;
    		:NO2DOAS.sigma.a4 = "0.015625" ;
    		:NO2DOAS.sigma.a5 = "0.015625" ;
    		:NO2DOAS.sigma.c0 = "1.0" ;
    		:NO2DOAS.sigma.c1 = "0.125" ;
    		:NO2DOAS.sigma.c2 = "0.015625" ;
    		:NO2DOAS.sigma.c3 = "0.015625" ;
    		:NO2DOAS.sigma.ring = "0.2" ;
    		:NO2DOAS.species = "NO2, O3, O2O2, H2O_vapor, H2O_liquid" ;
    		:NO2DOAS.wavelength_end = "465.0" ;
    		:NO2DOAS.wavelength_start = "405.0" ;
    		:NO2DOAS.write_diagnostic_output = "true" ;
    		:configuration.version.algorithm = "1.6.0" ;
    		:configuration.version.framework = "1.2.0" ;
    		:input.1.band = "4" ;
    		:input.1.irrType = "L1B_IR_UVN" ;
    		:input.1.type = "L1B_RA_BD4" ;
    		:input.2.band = "6" ;
    		:input.2.required = "false" ;
    		:input.2.type = "L2__FRESCO" ;
    		:input.3.band = "3" ;
    		:input.3.type = "L2__AER_AI" ;
    		:input.4.band = "3" ;
    		:input.4.required = "false" ;
    		:input.4.type = "L2__CLOUD_" ;
    		:input.5.band = "4" ;
    		:input.5.required = "false" ;
    		:input.5.type = "L2__O22CLD" ;
    		:input.count = "5" ;
    		:output.1.band = "4" ;
    		:output.1.config = "cfg/product/product.NO2O22.xml" ;
    		:output.1.level = "0" ;
    		:output.1.type = "L2__NO2___" ;
    		:output.compressionLevel = "3" ;
    		:output.count = "1" ;
    		:output.histogram.nitrogendioxide_stratospheric_column.logarithmic = "false" ;
    		:output.histogram.nitrogendioxide_stratospheric_column.range = "0,0.000166054" ;
    		:output.histogram.nitrogendioxide_total_column.logarithmic = "true" ;
    		:output.histogram.nitrogendioxide_total_column.range = "1.66054e-06,0.00166054" ;
    		:output.histogram.nitrogendioxide_tropospheric_column.logarithmic = "true" ;
    		:output.histogram.nitrogendioxide_tropospheric_column.range = "1.66054e-06,0.00166054" ;
    		:output.useCompression = "true" ;
    		:output.useFletcher32 = "true" ;
    		:output.useShuffleFilter = "true" ;
    		:processing.NO2_scd_limit = "-20.0e-6" ;
    		:processing.albedo_wavelength = "440.0" ;
    		:processing.albedo_wavelength_o2o2 = "475.0" ;
    		:processing.albedo_wavelengths = "463.0, 494.0" ;
    		:processing.algorithm = "NO2___" ;
    		:processing.cloud_selection = "0" ;
    		:processing.cloud_wavelength = "440.0" ;
    		:processing.cloud_wavelength_delta = "1.0" ;
    		:processing.correct_surface_pressure_for_altitude = "true" ;
    		:processing.dler.fractional_snice = "false" ;
    		:processing.dler.ice_max_threshold = "1" ;
    		:processing.dler.snow_max_threshold = "10" ;
    		:processing.dler.spatial_interpolation = "true" ;
    		:processing.dler.useDLER = "true" ;
    		:processing.dler.wavelengths = "440, 463, 494" ;
    		:processing.fitWindowExtent = "3" ;
    		:processing.groupDem = "DEM_RADIUS_05000" ;
    		:processing.irradFluxVarName = "irradiance_flux_cf" ;
    		:processing.radRingFluxVarName = "radiance_ring_flux_cf" ;
    		:processing.radianceFractionMinError = "0.4" ;
    		:processing.radianceFractionMinWarning = "0.8" ;
    		:processing.reflectance_from_model = "true" ;
    		:processing.reflectance_noise_floor = "2500.0" ;
    		:processing.saturationMaxFraction = "0.25" ;
    		:processing.saturationMaxWarningFraction = "0.0" ;
    		:processing.szaMax = "88.0" ;
    		:processing.szaMin = "0.0" ;
    		:processing.use_error_in_l1b = "false" ;
    		:processing.use_o22cld = "true" ;
    		:processing.use_spline_for_mu0 = "false" ;
    		:processing.vzaMax = "75.0" ;
    		:processing.vzaMin = "0.0" ;
    		:qa_value.AAI_warning = "100.0" ;
    		:qa_value.altitude_consistency_warning = "100.0" ;
    		:qa_value.amf_trop_geo_ratio_modification_percent = "45.0" ;
    		:qa_value.amf_trop_geo_ratio_threshold = "0.1" ;
    		:qa_value.cloud_radiance_fraction_modification_percent = "74.0" ;
    		:qa_value.cloud_radiance_fraction_threshold = "0.5" ;
    		:qa_value.cloud_warning = "100.0" ;
    		:qa_value.data_range_warning = "100.0" ;
    		:qa_value.deconvolution_warning = "100.0" ;
    		:qa_value.extrapolation_warning = "100.0" ;
    		:qa_value.input_spectrum_warning = "100.0" ;
    		:qa_value.interpolation_warning = "90.0" ;
    		:qa_value.low_cloud_fraction_warning = "100.0" ;
    		:qa_value.maximum_aerosol_index_modification_percent = "40.0" ;
    		:qa_value.maximum_aerosol_index_threshold = "1.0e10" ;
    		:qa_value.minimum_scene_pressure_modification_percent = "25.0" ;
    		:qa_value.minimum_scene_pressure_threshold = "30000.0" ;
    		:qa_value.no2_scd_precision_modification_percent = "15.0" ;
    		:qa_value.no2_scd_precision_threshold = "33.0e-6" ;
    		:qa_value.pixel_level_input_data_missing = "90.0" ;
    		:qa_value.signal_to_noise_ratio_warning = "100.0" ;
    		:qa_value.snow_ice_max_modification_percent = "73.0" ;
    		:qa_value.snow_ice_max_threshold = "1" ;
    		:qa_value.snow_ice_nocloud_modification_percent = "88" ;
    		:qa_value.snow_ice_nocloud_scene_pressure_fraction_threshold = "0.96" ;
    		:qa_value.snow_ice_nocloud_snow_threshold = "80" ;
    		:qa_value.snow_ice_warning = "100.0" ;
    		:qa_value.so2_volcanic_origin_certain_warning = "100.0" ;
    		:qa_value.so2_volcanic_origin_likely_warning = "100.0" ;
    		:qa_value.south_atlantic_anomaly_warning = "95.0" ;
    		:qa_value.sun_glint_correction = "100.0" ;
    		:qa_value.sun_glint_warning = "93.0" ;
    		:qa_value.surface_albedo_modification_percent = "20.0" ;
    		:qa_value.surface_albedo_threshold = "0.3" ;
    		:qa_value.sza_max_1_modification_percent = "30.0" ;
    		:qa_value.sza_max_1_threshold = "81.2" ;
    		:qa_value.sza_max_2_modification_percent = "10.0" ;
    		:qa_value.sza_max_2_threshold = "84.5" ;
    		:qa_value.thermal_instability_warning = "100.0" ;
    		:qa_value.wavelength_calibration_warning = "100.0" ;
    		:quality_control.missing_input.max_fraction = "0.25" ;
    		:quality_control.missing_scanlines.max_count = "60" ;
    		:quality_control.missing_scanlines.max_fraction = "0.05" ;
    		:quality_control.qa_value.limit = "0.5" ;
    		:quality_control.success.min_fraction = "0.001" ;
    		:wavelength_calibration.convergence_threshold = "1.0" ;
    		:wavelength_calibration.include_ring = "yes" ;
    		:wavelength_calibration.include_stretch = "no" ;
    		:wavelength_calibration.initial_guess.a0 = "1.0" ;
    		:wavelength_calibration.initial_guess.a1 = "0.1" ;
    		:wavelength_calibration.initial_guess.a2 = "0.01" ;
    		:wavelength_calibration.initial_guess.ring = "0.06" ;
    		:wavelength_calibration.initial_guess.shift = "0.0" ;
    		:wavelength_calibration.initial_guess.stretch = "0.0" ;
    		:wavelength_calibration.irr.include_ring = "no" ;
    		:wavelength_calibration.max_iterations = "12" ;
    		:wavelength_calibration.perform_wavelength_fit = "yes" ;
    		:wavelength_calibration.polynomial_order = "2" ;
    		:wavelength_calibration.sigma.a0 = "1.0" ;
    		:wavelength_calibration.sigma.a1 = "0.1" ;
    		:wavelength_calibration.sigma.a2 = "0.01" ;
    		:wavelength_calibration.sigma.ring = "0.06" ;
    		:wavelength_calibration.sigma.shift = "0.07" ;
    		:wavelength_calibration.sigma.stretch = "0.07" ;
    		:wavelength_calibration.window = "405.0, 465.0" ;
    		:wavelength_calibration_o22cld.convergence_threshold = "1.0" ;
    		:wavelength_calibration_o22cld.include_ring = "yes" ;
    		:wavelength_calibration_o22cld.include_stretch = "no" ;
    		:wavelength_calibration_o22cld.initial_guess.a0 = "1.0" ;
    		:wavelength_calibration_o22cld.initial_guess.a1 = "0.1" ;
    		:wavelength_calibration_o22cld.initial_guess.a2 = "0.01" ;
    		:wavelength_calibration_o22cld.initial_guess.ring = "0.06" ;
    		:wavelength_calibration_o22cld.initial_guess.shift = "0.0" ;
    		:wavelength_calibration_o22cld.initial_guess.stretch = "0.0" ;
    		:wavelength_calibration_o22cld.irr.include_ring = "no" ;
    		:wavelength_calibration_o22cld.max_iterations = "12" ;
    		:wavelength_calibration_o22cld.perform_wavelength_fit = "yes" ;
    		:wavelength_calibration_o22cld.polynomial_order = "2" ;
    		:wavelength_calibration_o22cld.sigma.a0 = "1.0" ;
    		:wavelength_calibration_o22cld.sigma.a1 = "0.1" ;
    		:wavelength_calibration_o22cld.sigma.a2 = "0.01" ;
    		:wavelength_calibration_o22cld.sigma.ring = "0.06" ;
    		:wavelength_calibration_o22cld.sigma.shift = "0.07" ;
    		:wavelength_calibration_o22cld.sigma.stretch = "0.07" ;
    		:wavelength_calibration_o22cld.window = "460.0, 490.0" ;
    		:joborder.processing.threads = "26" ;
    } // group ALGORITHM_SETTINGS

  group: GRANULE_DESCRIPTION {

    // group attributes:
    		:GranuleStart = "2024-01-24T06:39:07Z" ;
    		:GranuleEnd = "2024-01-24T06:44:18Z" ;
    		:InstrumentName = "TROPOMI" ;
    		:MissionName = "Sentinel-5 precursor" ;
    		:MissionShortName = "S5P" ;
    		:ProcessLevel = "2" ;
    		:ProcessingCenter = "PDGS-OP" ;
    		:ProcessingNode = "s5p-ops2-nrt-pn04" ;
    		:ProcessorVersion = "2.6.0" ;
    		:ProductFormatVersion = 20400 ;
    		:ProcessingMode = "Near-realtime" ;
    		:LongitudeOfDaysideNadirEquatorCrossing = 9.96921e+36f ;
    		:CollectionIdentifier = "03" ;
    		:ProductShortName = "L2__NO2___" ;
    } // group GRANULE_DESCRIPTION

  group: ISO_METADATA {

    // group attributes:
    		:gmd\:dateStamp = "2015-10-16" ;
    		:gmd\:fileIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__NO2___" ;
    		:gmd\:hierarchyLevelName = "EO Product Collection" ;
    		:gmd\:metadataStandardName = "ISO 19115-2 Geographic Information - Metadata Part 2 Extensions for imagery and gridded data" ;
    		:gmd\:metadataStandardVersion = "ISO 19115-2:2009(E), S5P profile" ;
    		:objectType = "gmi:MI_Metadata" ;

    group: gmd\:language {

      // group attributes:
      		:codeList = "http://www.loc.gov/standards/iso639-2/" ;
      		:codeListValue = "eng" ;
      		:objectType = "gmd:LanguageCode" ;
      } // group gmd\:language

    group: gmd\:characterSet {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
      		:codeListValue = "utf8" ;
      		:objectType = "gmd:MD_CharacterSetCode" ;
      } // group gmd\:characterSet

    group: gmd\:hierarchyLevel {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
      		:codeListValue = "series" ;
      		:objectType = "gmd:MD_ScopeCode" ;
      } // group gmd\:hierarchyLevel

    group: gmd\:contact {

      // group attributes:
      		:gmd\:organisationName = "Copernicus Space Component Data Access System,  ESA, Services Coordinated Interface" ;
      		:objectType = "gmd:CI_ResponsibleParty" ;

      group: gmd\:contactInfo {

        // group attributes:
        		:objectType = "gmd:CI_Contact" ;

        group: gmd\:address {

          // group attributes:
          		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
          		:objectType = "gmd:CI_Address" ;
          } // group gmd\:address
        } // group gmd\:contactInfo

      group: gmd\:role {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
        		:codeListValue = "pointOfContact" ;
        		:objectType = "gmd:CI_RoleCode" ;
        } // group gmd\:role
      } // group gmd\:contact

    group: gmd\:identificationInfo {

      // group attributes:
      		:gmd\:abstract = "Nitrogen dioxide tropospheric column with a spatial resolution of 5.5x3.5 km2 observed at about 13:30 local solar time from spectra measured by TROPOMI" ;
      		:gmd\:credit = "The Sentinel 5 Precursor TROPOMI Level 2 products are developed with funding from the European Space Agency (ESA), the Netherlands Space Office (NSO), the Belgian Science Policy Office, the German Aerospace Center (DLR) and the Bayerisches Staatsministerium für Wirtschaft und Medien, Energie und Technologie (StMWi)." ;
      		:gmd\:language = "eng" ;
      		:gmd\:topicCategory = "climatologyMeteorologyAtmosphere" ;
      		:objectType = "gmd:MD_DataIdentification" ;

      group: gmd\:citation {

        // group attributes:
        		:gmd\:title = "TROPOMI/S5P NO2 5-minute L2 Swath 5.5x3.5km" ;
        		:objectType = "gmd:CI_Citation" ;

        group: gmd\:date {

          // group attributes:
          		:gmd\:date = "2024-01-24" ;
          		:objectType = "gmd:CI_Date" ;

          group: gmd\:dateType {

            // group attributes:
            		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
            		:codeListValue = "creation" ;
            		:objectType = "gmd:CI_DateTypeCode" ;
            } // group gmd\:dateType
          } // group gmd\:date

        group: gmd\:identifier {

          // group attributes:
          		:gmd\:code = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__NO2___" ;
          		:objectType = "gmd:MD_Identifier" ;
          } // group gmd\:identifier
        } // group gmd\:citation

      group: gmd\:pointOfContact {

        // group attributes:
        		:gmd\:organisationName = "Copernicus Space Component Data Access System,  ESA, Services Coordinated Interface" ;
        		:objectType = "gmd:CI_ResponsibleParty" ;

        group: gmd\:contactInfo {

          // group attributes:
          		:objectType = "gmd:CI_Contact" ;

          group: gmd\:address {

            // group attributes:
            		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
            		:objectType = "gmd:CI_Address" ;
            } // group gmd\:address
          } // group gmd\:contactInfo

        group: gmd\:role {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
          		:codeListValue = "distributor" ;
          		:objectType = "gmd:CI_RoleCode" ;
          } // group gmd\:role
        } // group gmd\:pointOfContact

      group: gmd\:descriptiveKeywords\#1 {

        // group attributes:
        		:gmd\:keyword\#1 = "Atmospheric conditions" ;
        		:objectType = "gmd:MD_Keywords" ;

        group: gmd\:type {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode" ;
          		:codeListValue = "theme" ;
          		:objectType = "gmd:MD_KeywordTypeCode" ;
          } // group gmd\:type

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "GEMET - INSPIRE themes, version 1.0" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2008-06-01" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName
        } // group gmd\:descriptiveKeywords\#1

      group: gmd\:descriptiveKeywords\#2 {

        // group attributes:
        		:gmd\:keyword\#1 = "troposphere_mole_content_of_nitrogen_dioxide" ;
        		:objectType = "gmd:MD_Keywords" ;
        		:gmd\:keyword\#2 = "stratosphere_mole_content_of_nitrogen_dioxide" ;
        		:gmd\:keyword\#3 = "atmosphere_mole_content_of_nitrogen_dioxide" ;

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "CF Standard Name Table v65" ;
          		:xlink\:href = "http://cfconventions.org/standard-names.html" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2019-04-09" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName
        } // group gmd\:descriptiveKeywords\#2

      group: gmd\:resourceConstraints {

        // group attributes:
        		:gmd\:useLimitation = "no conditions apply" ;
        		:objectType = "gmd:MD_LegalConstraints" ;

        group: gmd\:accessConstraints {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_RestrictionCode" ;
          		:codeListValue = "copyright" ;
          		:objectType = "gmd:MD_RestrictionCode" ;
          } // group gmd\:accessConstraints
        } // group gmd\:resourceConstraints

      group: gmd\:spatialRepresentationType {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_SpatialRepresentationTypeCode" ;
        		:codeListValue = "grid" ;
        		:objectType = "gmd:MD_SpatialRepresentationTypeCode" ;
        } // group gmd\:spatialRepresentationType

      group: gmd\:characterSet {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
        		:codeListValue = "utf8" ;
        		:objectType = "gmd:MD_CharacterSetCode" ;
        } // group gmd\:characterSet

      group: gmd\:extent {

        // group attributes:
        		:objectType = "gmd:EX_Extent" ;

        group: gmd\:geographicElement {

          // group attributes:
          		:gmd\:eastBoundLongitude = 111.3999f ;
          		:gmd\:northBoundLatitude = 56.08662f ;
          		:gmd\:southBoundLatitude = 32.02938f ;
          		:gmd\:westBoundLongitude = 71.52991f ;
          		:gmd\:extentTypeCode = "true" ;
          		:objectType = "gmd:EX_GeographicBoundingBox" ;
          } // group gmd\:geographicElement

        group: gmd\:temporalElement {

          // group attributes:
          		:objectType = "gmd:EX_TemporalExtent" ;

          group: gmd\:extent {

            // group attributes:
            		:gml\:beginPosition = "2024-01-24T06:39:07Z" ;
            		:gml\:endPosition = "2024-01-24T06:44:18Z" ;
            		:objectType = "gml:TimePeriod" ;
            } // group gmd\:extent
          } // group gmd\:temporalElement
        } // group gmd\:extent
      } // group gmd\:identificationInfo

    group: gmd\:dataQualityInfo {

      // group attributes:
      		:objectType = "gmd:DQ_DataQuality" ;

      group: gmd\:scope {

        // group attributes:
        		:objectType = "gmd:DQ_Scope" ;

        group: gmd\:level {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
          		:codeListValue = "dataset" ;
          		:objectType = "gmd:MD_ScopeCode" ;
          } // group gmd\:level
        } // group gmd\:scope

      group: gmd\:report {

        // group attributes:
        		:objectType = "gmd:DQ_DomainConsistency" ;

        group: gmd\:result {

          // group attributes:
          		:objectType = "gmd:DQ_ConformanceResult" ;
          		:gmd\:pass = "true" ;
          		:gmd\:explanation = "INSPIRE Data specification for orthoimagery is not yet officially published so conformity has not yet been evaluated" ;

          group: gmd\:specification {

            // group attributes:
            		:objectType = "gmd:CI_Citation" ;
            		:gmd\:title = "INSPIRE Data Specification on Orthoimagery - Guidelines, version 3.0rc3" ;

            group: gmd\:date {

              // group attributes:
              		:gmd\:date = "2013-02-04" ;
              		:objectType = "gmd:CI_Date" ;

              group: gmd\:dateType {

                // group attributes:
                		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                		:codeListValue = "publication" ;
                		:objectType = "gmd:CI_DateTypeCode" ;
                } // group gmd\:dateType
              } // group gmd\:date
            } // group gmd\:specification
          } // group gmd\:result
        } // group gmd\:report

      group: gmd\:lineage {

        // group attributes:
        		:objectType = "gmd:LI_Lineage" ;
        		:gmd\:statement = "L2 NO2___ dataset produced by PDGS-OP from the S5P/TROPOMI L1B product" ;

        group: gmd\:processStep {

          // group attributes:
          		:objectType = "gmi:LE_ProcessStep" ;
          		:gmd\:description = "Processing of L1b to L2 NO2___ data for orbit 32544 using the KNMI processor version 2.6.0" ;

          group: gmi\:output {

            // group attributes:
            		:gmd\:description = "TROPOMI/S5P NO2 5-minute L2 Swath 5.5x3.5km" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmd\:sourceCitation {

              // group attributes:
              		:gmd\:title = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24" ;
                		:objectType = "gmd:CI_DateTime" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:identifier {

                // group attributes:
                		:gmd\:code = "L2__NO2___" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmd\:identifier
              } // group gmd\:sourceCitation

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L2" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel
            } // group gmi\:output

          group: gmi\:processingInformation {

            // group attributes:
            		:objectType = "gmi:LE_Processing" ;

            group: gmi\:identifier {

              // group attributes:
              		:gmd\:code = "KNMI L2 NO2___ processor, version 2.6.0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:identifier

            group: gmi\:softwareReference {

              // group attributes:
              		:gmd\:title = "TROPNLL2DP processor" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2023-09-28T07:04:00Z" ;
                		:objectType = "gmd:CI_DateTime" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:softwareReference

            group: gmi\:documentation\#1 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "TROPOMI ATBD of the total and tropospheric NO2 data products; S5P-KNMI-L2-0005-RP; release 1.0" ;
              		:doi = "N/A" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-30" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "revision" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#1

            group: gmi\:documentation\#2 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual Nitrogen Dioxide; S5P-KNMI-L2-0021-MA; release 1.0" ;
              		:doi = "N/A" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-30" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "revision" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#2
            } // group gmi\:processingInformation

          group: gmi\:report {

            // group attributes:
            		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the KNMI L2 NO2___ processor" ;
            		:gmi\:fileType = "netCDF-4" ;
            		:gmi\:name = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919.nc" ;
            		:objectType = "gmi:LE_ProcessStepReport" ;
            } // group gmi\:report

          group: gmd\:source\#1 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary CTM AUX_CTMFCT model input data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary CTM AUX_CTMFCT model input data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_AUX_CTMFCT_20240124T000000_20240125T000000_20240124T060507.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#1

          group: gmd\:source\#2 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L4" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20240124T030000_20240124T120000_20240124T000000.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#2

          group: gmd\:source\#3 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L4" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_TP_20240124T030000_20240124T120000_20240124T000000.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#3

          group: gmd\:source\#4 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary AUX_O3___M reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary AUX_O3___M reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_AUX_O3___M_00000000T000000_99999999T999999_20210119T232003.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#4

          group: gmd\:source\#5 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Processor CFG_NO2___ configuration file" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Processor CFG_NO2___ configuration file" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_CFG_NO2____00000000T000000_99999999T999999_20230901T000000.cfg" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#5

          group: gmd\:source\#6 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_IR_UVN_20240123T105621_20240123T123751_32533_03_020100_20240123T142235.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#6

          group: gmd\:source\#7 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD4 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD4 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD4_20240124T063906_20240124T064418_32544_03_020100_20240124T065843.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#7

          group: gmd\:source\#8 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__AER_AI product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__AER_AI product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L2__AER_AI_20240124T063912_20240124T064412_32544_03_020600_20240124T071559.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#8

          group: gmd\:source\#9 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__FRESCO product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__FRESCO product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L2__FRESCO_20240124T063912_20240124T064412_32544_03_020600_20240124T071554.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#9

          group: gmd\:source\#10 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary LUT_NO2AMF algorithm lookup table" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary LUT_NO2AMF algorithm lookup table" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_LUT_NO2AMF_00000000T000000_99999999T999999_20160527T173500.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#10

          group: gmd\:source\#11 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary LUT_NO2CLD algorithm lookup table" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary LUT_NO2CLD algorithm lookup table" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_LUT_NO2CLD_00000000T000000_99999999T999999_20191115T193538.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#11

          group: gmd\:source\#12 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary LUT_O22CLD algorithm lookup table" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary LUT_O22CLD algorithm lookup table" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_LUT_O22CLD_00000000T000000_99999999T999999_20200305T174212.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#12

          group: gmd\:source\#13 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_DEM___ reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_DEM___ reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_DEM____20190404T150000_99999999T999999_20190405T143622.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#13

          group: gmd\:source\#14 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_LER___ reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_LER___ reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_LER____00000000T000000_99999999T999999_20220113T000000.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#14

          group: gmd\:source\#15 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_SOLAR_ reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_SOLAR_ reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_SOLAR__00000000T000000_99999999T999999_20210107T132455.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#15

          group: gmd\:source\#16 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_XS_NO2 reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-01-24T07:22:46Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_XS_NO2 reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_XS_NO2_00000000T000000_99999999T999999_20180118T134308.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#16
          } // group gmd\:processStep
        } // group gmd\:lineage
      } // group gmd\:dataQualityInfo

    group: gmi\:acquisitionInformation {

      // group attributes:
      		:objectType = "gmi:MI_AcquisitionInformation" ;

      group: gmi\:platform {

        // group attributes:
        		:gmi\:description = "Sentinel 5 Precursor" ;
        		:objectType = "gmi:MI_Platform" ;

        group: gmi\:identifier {

          // group attributes:
          		:gmd\:code = "S5P" ;
          		:gmd\:codeSpace = "http://www.esa.int/" ;
          		:objectType = "gmd:RS_Identifier" ;
          } // group gmi\:identifier

        group: gmi\:instrument {

          // group attributes:
          		:objectType = "gmi:MI_Instrument" ;
          		:gmi\:type = "UV-VIS-NIR-SWIR imaging spectrometer" ;

          group: gmi\:identifier {

            // group attributes:
            		:gmd\:code = "TROPOMI" ;
            		:gmd\:codeSpace = "http://www.esa.int/" ;
            		:objectType = "gmd:RS_Identifier" ;
            } // group gmi\:identifier
          } // group gmi\:instrument
        } // group gmi\:platform
      } // group gmi\:acquisitionInformation
    } // group ISO_METADATA

  group: EOP_METADATA {

    // group attributes:
    		:gml\:id = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919.ID" ;
    		:objectType = "atm:EarthObservation" ;

    group: om\:phenomenonTime {

      // group attributes:
      		:gml\:beginPosition = "2024-01-24T06:39:07Z" ;
      		:gml\:endPosition = "2024-01-24T06:44:18Z" ;
      		:objectType = "gml:TimePeriod" ;
      } // group om\:phenomenonTime

    group: om\:procedure {

      // group attributes:
      		:gml\:id = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919.EOE" ;
      		:objectType = "eop:EarthObservationEquipment" ;

      group: eop\:platform {

        // group attributes:
        		:eop\:shortName = "Sentinel-5p" ;
        		:objectType = "eop:Platform" ;
        } // group eop\:platform

      group: eop\:instrument {

        // group attributes:
        		:eop\:shortName = "TROPOMI" ;
        		:objectType = "eop:Instrument" ;
        } // group eop\:instrument

      group: eop\:sensor {

        // group attributes:
        		:eop\:sensorType = "ATMOSPHERIC" ;
        		:objectType = "eop:Sensor" ;
        } // group eop\:sensor

      group: eop\:acquisitionParameters {

        // group attributes:
        		:eop\:orbitNumber = 32544 ;
        		:objectType = "eop:Acquisition" ;
        } // group eop\:acquisitionParameters
      } // group om\:procedure

    group: om\:observedProperty {

      // group attributes:
      		:nilReason = "inapplicable" ;
      } // group om\:observedProperty

    group: om\:featureOfInterest {

      // group attributes:
      		:objectType = "eop:FootPrint" ;
      		:gml\:id = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919.FP" ;

      group: eop\:multiExtentOf {

        // group attributes:
        		:objectType = "gml:MultiSurface" ;

        group: gml\:surfaceMembers {

          // group attributes:
          		:objectType = "gml:Polygon" ;

          group: gml\:exterior {

            // group attributes:
            		:gml\:posList = "48.783443 71.529915 47.488457 72.689064 46.18085 73.78759 44.86121 74.82913 43.530632 75.81823 42.19012 76.75907 40.840424 77.65491 39.482502 78.50974 38.116737 79.3258 36.74376 80.105835 35.364304 80.852745 33.97872 81.56859 32.587418 82.25546 32.029385 82.52248 32.072224 82.60929 32.84438 84.21279 34.040558 86.87922 34.74118 88.59043 35.328728 90.157455 35.726097 91.31642 36.09224 92.48481 36.3584 93.41609 36.618156 94.41427 36.8164 95.25397 37.001934 96.12058 37.017853 96.199356 37.176773 97.03294 37.34222 98.01611 37.474583 98.92516 37.61231 100.05274 37.72015 101.15417 37.825672 102.60944 37.896538 104.14198 37.937424 106.37593 37.905827 109.07682 37.819588 111.39986 39.26621 111.2492 40.71214 111.106834 42.15733 110.97393 43.60175 110.850334 45.04542 110.737045 46.488308 110.634705 47.930305 110.544266 49.371513 110.46658 50.811737 110.40257 52.251087 110.353714 53.689312 110.32182 55.126568 110.30872 55.70121 110.30876 55.71321 110.16405 55.91502 107.266365 56.07449 102.922874 56.078316 100.168755 56.00846 97.690895 55.909184 95.89492 55.766857 94.122246 55.62285 92.73961 55.438763 91.28952 55.26065 90.09612 55.055225 88.890305 55.03549 88.782005 54.816 87.64944 54.532757 86.34513 54.248222 85.16925 53.86642 83.750046 53.46436 82.40421 52.89251 80.683365 52.245213 78.93529 51.22892 76.48924 49.898735 73.66475 48.783443 71.529915 48.783443 71.529915" ;
            		:objectType = "gml:LinearRing" ;
            } // group gml\:exterior
          } // group gml\:surfaceMembers
        } // group eop\:multiExtentOf
      } // group om\:featureOfInterest

    group: eop\:metaDataProperty {

      // group attributes:
      		:objectType = "eop:EarthObservationMetaData" ;
      		:eop\:acquisitionType = "NOMINAL" ;
      		:eop\:identifier = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919" ;
      		:eop\:doi = "N/A" ;
      		:eop\:parentIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__NO2___" ;
      		:eop\:productType = "S5P_NRTI_NO2___" ;
      		:eop\:status = "ACQUIRED" ;
      		:eop\:productQualityStatus = "NOMINAL" ;
      		:eop\:productQualityDegradationTag = "NOT APPLICABLE" ;

      group: eop\:processing {

        // group attributes:
        		:objectType = "eop:ProcessingInformation" ;
        		:eop\:processingCenter = "PDGS-OP" ;
        		:eop\:processingDate = "2024-01-24" ;
        		:eop\:processingLevel = "L2" ;
        		:eop\:processorName = "TROPNLL2DP" ;
        		:eop\:processorVersion = "2.6.0" ;
        		:eop\:nativeProductFormat = "netCDF-4" ;
        		:eop\:processingMode = "NRTI" ;
        } // group eop\:processing
      } // group eop\:metaDataProperty
    } // group EOP_METADATA

  group: ESA_METADATA {

    group: earth_explorer_header {

      // group attributes:
      		:objectType = "Earth_Explorer_Header" ;

      group: fixed_header {

        // group attributes:
        		:objectType = "Fixed_Header" ;
        		:File_Name = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919" ;
        		:File_Description = "Nitrogen dioxide tropospheric column with a spatial resolution of 5.5x3.5 km2 observed at about 13:30 local solar time from spectra measured by TROPOMI" ;
        		:Notes = "" ;
        		:Mission = "S5P" ;
        		:File_Class = "NRTI" ;
        		:File_Type = "L2__NO2___" ;
        		:File_Version = 1 ;

        group: validity_period {

          // group attributes:
          		:objectType = "Validity_Period" ;
          		:Validity_Start = "UTC=2024-01-24T06:39:07" ;
          		:Validity_Stop = "UTC=2024-01-24T06:44:18" ;
          } // group validity_period

        group: source {

          // group attributes:
          		:objectType = "Source" ;
          		:System = "PDGS-OP" ;
          		:Creator = "TROPNLL2DP" ;
          		:Creator_Version = "2.6.0" ;
          		:Creation_Date = "UTC=2024-01-24T07:20:29" ;
          } // group source
        } // group fixed_header

      group: variable_header {

        // group attributes:
        		:objectType = "Variable_Header" ;

        group: gmd\:lineage {

          // group attributes:
          		:objectType = "gmd:LI_Lineage" ;
          		:gmd\:statement = "L2 NO2___ dataset produced by PDGS-OP from the S5P/TROPOMI L1B product" ;

          group: gmd\:processStep {

            // group attributes:
            		:objectType = "gmi:LE_ProcessStep" ;
            		:gmd\:description = "Processing of L1b to L2 NO2___ data for orbit 32544 using the KNMI processor version 2.6.0" ;

            group: gmi\:output {

              // group attributes:
              		:gmd\:description = "TROPOMI/S5P NO2 5-minute L2 Swath 5.5x3.5km" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmd\:sourceCitation {

                // group attributes:
                		:gmd\:title = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:identifier {

                  // group attributes:
                  		:gmd\:code = "L2__NO2___" ;
                  		:objectType = "gmd:MD_Identifier" ;
                  } // group gmd\:identifier
                } // group gmd\:sourceCitation

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L2" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel
              } // group gmi\:output

            group: gmi\:processingInformation {

              // group attributes:
              		:objectType = "gmi:LE_Processing" ;

              group: gmi\:identifier {

                // group attributes:
                		:gmd\:code = "KNMI L2 NO2___ processor, version 2.6.0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:identifier

              group: gmi\:softwareReference {

                // group attributes:
                		:gmd\:title = "TROPNLL2DP processor" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2023-09-28T07:04:00Z" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:softwareReference

              group: gmi\:documentation\#1 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "TROPOMI ATBD of the total and tropospheric NO2 data products; S5P-KNMI-L2-0005-RP; release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-30" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "revision" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#1

              group: gmi\:documentation\#2 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual Nitrogen Dioxide; S5P-KNMI-L2-0021-MA; release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-30" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "revision" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#2
              } // group gmi\:processingInformation

            group: gmi\:report {

              // group attributes:
              		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the KNMI L2 NO2___ processor" ;
              		:gmi\:fileType = "netCDF-4" ;
              		:gmi\:name = "S5P_NRTI_L2__NO2____20240124T063912_20240124T064412_32544_03_020600_20240124T071919.nc" ;
              		:objectType = "gmi:LE_ProcessStepReport" ;
              } // group gmi\:report

            group: gmd\:source\#1 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary CTM AUX_CTMFCT model input data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary CTM AUX_CTMFCT model input data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_CTMFCT_20240124T000000_20240125T000000_20240124T060507.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#1

            group: gmd\:source\#2 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L4" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20240124T030000_20240124T120000_20240124T000000.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#2

            group: gmd\:source\#3 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L4" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_TP_20240124T030000_20240124T120000_20240124T000000.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#3

            group: gmd\:source\#4 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary AUX_O3___M reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary AUX_O3___M reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_O3___M_00000000T000000_99999999T999999_20210119T232003.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#4

            group: gmd\:source\#5 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Processor CFG_NO2___ configuration file" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Processor CFG_NO2___ configuration file" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_CFG_NO2____00000000T000000_99999999T999999_20230901T000000.cfg" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#5

            group: gmd\:source\#6 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_IR_UVN_20240123T105621_20240123T123751_32533_03_020100_20240123T142235.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#6

            group: gmd\:source\#7 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD4 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD4 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD4_20240124T063906_20240124T064418_32544_03_020100_20240124T065843.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#7

            group: gmd\:source\#8 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__AER_AI product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__AER_AI product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L2__AER_AI_20240124T063912_20240124T064412_32544_03_020600_20240124T071559.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#8

            group: gmd\:source\#9 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__FRESCO product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__FRESCO product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L2__FRESCO_20240124T063912_20240124T064412_32544_03_020600_20240124T071554.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#9

            group: gmd\:source\#10 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_NO2AMF algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_NO2AMF algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_NO2AMF_00000000T000000_99999999T999999_20160527T173500.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#10

            group: gmd\:source\#11 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_NO2CLD algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_NO2CLD algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_NO2CLD_00000000T000000_99999999T999999_20191115T193538.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#11

            group: gmd\:source\#12 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_O22CLD algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_O22CLD algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_O22CLD_00000000T000000_99999999T999999_20200305T174212.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#12

            group: gmd\:source\#13 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_DEM___ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_DEM___ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_DEM____20190404T150000_99999999T999999_20190405T143622.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#13

            group: gmd\:source\#14 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_LER___ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_LER___ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_LER____00000000T000000_99999999T999999_20220113T000000.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#14

            group: gmd\:source\#15 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_SOLAR_ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_SOLAR_ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_SOLAR__00000000T000000_99999999T999999_20210107T132455.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#15

            group: gmd\:source\#16 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_XS_NO2 reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-01-24T07:22:46Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_XS_NO2 reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_XS_NO2_00000000T000000_99999999T999999_20180118T134308.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#16
            } // group gmd\:processStep
          } // group gmd\:lineage

        group: subsystem_information {

          // group attributes:
          		:objectType = "subsystem_information" ;

          group: subsystem\#0 {

            // group attributes:
            		:Authors = "H.J. Eskes, K.F. Boersma, J.D. Maasakkers" ;
            		:Email = "eskes@knmi.nl" ;
            		:Institution = "KNMI (Royal Netherlands Meteorological Institute)" ;
            		:Name = "TM5-MP-Domino3" ;
            		:Version = "3.5.4" ;
            		:VersionDate = "2019-01-18" ;
            } // group subsystem\#0
          } // group subsystem_information
        } // group variable_header
      } // group earth_explorer_header
    } // group ESA_METADATA
  } // group METADATA
}
